`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Created for Indiana University's E315 Class
//
// 
// Andrew Lukefahr
// lukefahr@iu.edu
//
// 2021-03-24
// 2020-04-27
//
//////////////////////////////////////////////////////////////////////////////////

module dot_80_40(

		// AXI4-Stream Interface
		input                           clk,
		input                           rst,

        // Incomming Matrix AXI4-Stream
		input [31:0]                    INPUT_AXIS_TDATA,
        input                           INPUT_AXIS_TLAST,
        input                           INPUT_AXIS_TVALID,
        output                          INPUT_AXIS_TREADY,
        
        // Outgoing Vector AXI4-Stream 		
		output [31:0]                   OUTPUT_AXIS_TDATA,
        output                          OUTPUT_AXIS_TLAST,
        output                          OUTPUT_AXIS_TVALID,
        input                           OUTPUT_AXIS_TREADY 

    );
    
// This is autogenerated. See ../vtests/dot_80_40/dot_80_40.py for details. 
localparam ROWS = 80;
localparam COLS = 40;

localparam logic [31:0] weights [0:ROWS-1] [0:COLS-1] = '{
  '{ 
    $shortrealtobits(0.45885798),$shortrealtobits(0.09269916),$shortrealtobits(0.47095236),$shortrealtobits(-0.27914006),
    $shortrealtobits(-0.4357709),$shortrealtobits(0.37904724),$shortrealtobits(-0.29015967),$shortrealtobits(0.48655275),
    $shortrealtobits(0.33570504),$shortrealtobits(-0.141348),$shortrealtobits(-0.16425659),$shortrealtobits(0.37424883),
    $shortrealtobits(0.12360277),$shortrealtobits(0.22448532),$shortrealtobits(-0.027763547),$shortrealtobits(0.012192721),
    $shortrealtobits(-0.25464702),$shortrealtobits(-0.03298609),$shortrealtobits(-0.25456968),$shortrealtobits(0.32051057),
    $shortrealtobits(-0.2859922),$shortrealtobits(-0.4034654),$shortrealtobits(-0.2586356),$shortrealtobits(0.39009368),
    $shortrealtobits(0.28853428),$shortrealtobits(0.2839936),$shortrealtobits(0.0937717),$shortrealtobits(-0.06045808),
    $shortrealtobits(0.3494113),$shortrealtobits(0.121588804),$shortrealtobits(0.21573931),$shortrealtobits(-0.44571322),
    $shortrealtobits(-0.2645882),$shortrealtobits(0.37002876),$shortrealtobits(-0.0763041),$shortrealtobits(-0.095477),
    $shortrealtobits(-0.32527575),$shortrealtobits(-0.09613615),$shortrealtobits(-0.34059972),$shortrealtobits(-0.14155692)
  },
  '{ 
    $shortrealtobits(0.058472313),$shortrealtobits(0.14750688),$shortrealtobits(0.16937777),$shortrealtobits(-0.5251201),
    $shortrealtobits(-0.2299765),$shortrealtobits(-0.24935059),$shortrealtobits(0.43774527),$shortrealtobits(-0.07214785),
    $shortrealtobits(-0.19901769),$shortrealtobits(0.3520499),$shortrealtobits(0.056439083),$shortrealtobits(0.21418582),
    $shortrealtobits(-0.31059694),$shortrealtobits(0.15499203),$shortrealtobits(-0.24822634),$shortrealtobits(0.38136253),
    $shortrealtobits(0.4253648),$shortrealtobits(0.42777315),$shortrealtobits(-0.27873072),$shortrealtobits(-0.16869819),
    $shortrealtobits(-0.13061513),$shortrealtobits(-0.34887335),$shortrealtobits(0.046889763),$shortrealtobits(-0.4784313),
    $shortrealtobits(0.29052544),$shortrealtobits(0.14805283),$shortrealtobits(0.5058073),$shortrealtobits(0.23925963),
    $shortrealtobits(0.57548004),$shortrealtobits(-0.33365896),$shortrealtobits(-0.35804406),$shortrealtobits(0.07740109),
    $shortrealtobits(0.558082),$shortrealtobits(0.3264367),$shortrealtobits(0.017206598),$shortrealtobits(0.38324153),
    $shortrealtobits(-0.044437665),$shortrealtobits(-0.2013156),$shortrealtobits(0.28911883),$shortrealtobits(0.48443142)
  },
  '{ 
    $shortrealtobits(0.48097116),$shortrealtobits(-0.20028183),$shortrealtobits(-0.055972178),$shortrealtobits(0.31016755),
    $shortrealtobits(0.07261986),$shortrealtobits(-0.08674763),$shortrealtobits(0.03729569),$shortrealtobits(0.07724701),
    $shortrealtobits(-0.0016563042),$shortrealtobits(0.2780921),$shortrealtobits(-0.09847667),$shortrealtobits(0.22420877),
    $shortrealtobits(-0.15187259),$shortrealtobits(-0.14109828),$shortrealtobits(-0.19528754),$shortrealtobits(0.12981188),
    $shortrealtobits(-0.28370583),$shortrealtobits(-0.13403037),$shortrealtobits(0.337566),$shortrealtobits(0.113240525),
    $shortrealtobits(0.07131668),$shortrealtobits(0.1617904),$shortrealtobits(-0.288494),$shortrealtobits(-0.45081896),
    $shortrealtobits(0.39297736),$shortrealtobits(-0.4678036),$shortrealtobits(-0.5343804),$shortrealtobits(0.14880238),
    $shortrealtobits(-0.7801203),$shortrealtobits(-0.3195786),$shortrealtobits(-0.4200931),$shortrealtobits(-0.36821407),
    $shortrealtobits(-0.4246308),$shortrealtobits(0.28391415),$shortrealtobits(-0.29421163),$shortrealtobits(-0.20614783),
    $shortrealtobits(0.41660562),$shortrealtobits(-0.26203525),$shortrealtobits(-0.26258394),$shortrealtobits(-0.21484596)
  },
  '{ 
    $shortrealtobits(0.16808861),$shortrealtobits(-0.047700785),$shortrealtobits(-0.30293432),$shortrealtobits(0.54289997),
    $shortrealtobits(0.22124673),$shortrealtobits(-0.35519302),$shortrealtobits(-0.0625691),$shortrealtobits(-0.41093418),
    $shortrealtobits(0.07981887),$shortrealtobits(-0.08063049),$shortrealtobits(-0.12886913),$shortrealtobits(0.35807544),
    $shortrealtobits(0.46791637),$shortrealtobits(-0.4518445),$shortrealtobits(-0.20119022),$shortrealtobits(-0.2569115),
    $shortrealtobits(-0.39230675),$shortrealtobits(0.04657054),$shortrealtobits(-0.29183844),$shortrealtobits(0.034059934),
    $shortrealtobits(0.10895447),$shortrealtobits(-0.20255671),$shortrealtobits(0.29505566),$shortrealtobits(0.5036012),
    $shortrealtobits(0.33886838),$shortrealtobits(-0.50621),$shortrealtobits(0.058435507),$shortrealtobits(0.32703844),
    $shortrealtobits(0.37767732),$shortrealtobits(-0.27103233),$shortrealtobits(0.23019953),$shortrealtobits(0.43297467),
    $shortrealtobits(-0.53505737),$shortrealtobits(-0.12748961),$shortrealtobits(-0.1639826),$shortrealtobits(0.47773147),
    $shortrealtobits(0.19141494),$shortrealtobits(0.067063875),$shortrealtobits(0.51009643),$shortrealtobits(0.28296015)
  },
  '{ 
    $shortrealtobits(0.2430795),$shortrealtobits(0.44792315),$shortrealtobits(0.763975),$shortrealtobits(-0.06965235),
    $shortrealtobits(0.9541131),$shortrealtobits(0.1915156),$shortrealtobits(-0.051478922),$shortrealtobits(0.24432373),
    $shortrealtobits(0.5864828),$shortrealtobits(-0.032127727),$shortrealtobits(0.5441346),$shortrealtobits(-0.17603497),
    $shortrealtobits(0.32119995),$shortrealtobits(-0.042057794),$shortrealtobits(-0.20371997),$shortrealtobits(-0.047382236),
    $shortrealtobits(0.28870398),$shortrealtobits(0.097245775),$shortrealtobits(0.2748548),$shortrealtobits(-0.022933053),
    $shortrealtobits(-0.08351384),$shortrealtobits(0.4086131),$shortrealtobits(0.12909675),$shortrealtobits(0.020897266),
    $shortrealtobits(-0.16898784),$shortrealtobits(0.1654829),$shortrealtobits(0.36030704),$shortrealtobits(-0.76528305),
    $shortrealtobits(0.06916957),$shortrealtobits(-0.07844596),$shortrealtobits(-0.30489895),$shortrealtobits(-1.0374317),
    $shortrealtobits(0.2178733),$shortrealtobits(-0.31467804),$shortrealtobits(-0.0871871),$shortrealtobits(0.23576728),
    $shortrealtobits(-0.6258584),$shortrealtobits(-0.36045298),$shortrealtobits(0.08648108),$shortrealtobits(-0.028165584)
  },
  '{ 
    $shortrealtobits(0.42643276),$shortrealtobits(0.32872787),$shortrealtobits(-0.2415185),$shortrealtobits(0.17189324),
    $shortrealtobits(0.56030595),$shortrealtobits(0.35585067),$shortrealtobits(0.19265907),$shortrealtobits(0.21311097),
    $shortrealtobits(0.046162486),$shortrealtobits(0.30274493),$shortrealtobits(-0.2486716),$shortrealtobits(-0.39269862),
    $shortrealtobits(0.030138435),$shortrealtobits(0.3894209),$shortrealtobits(-0.19392566),$shortrealtobits(0.29585207),
    $shortrealtobits(-0.090557314),$shortrealtobits(-0.2535402),$shortrealtobits(0.14259475),$shortrealtobits(0.47398064),
    $shortrealtobits(0.03997285),$shortrealtobits(0.110087596),$shortrealtobits(0.46159816),$shortrealtobits(0.40776923),
    $shortrealtobits(0.49332365),$shortrealtobits(0.17731488),$shortrealtobits(0.46424335),$shortrealtobits(-0.16404793),
    $shortrealtobits(0.72305614),$shortrealtobits(0.39767665),$shortrealtobits(-0.555848),$shortrealtobits(0.26052985),
    $shortrealtobits(0.15525635),$shortrealtobits(-0.010110608),$shortrealtobits(-0.7336198),$shortrealtobits(0.20845065),
    $shortrealtobits(0.22280526),$shortrealtobits(-0.35965148),$shortrealtobits(-0.0127329),$shortrealtobits(0.0035724102)
  },
  '{ 
    $shortrealtobits(0.7090308),$shortrealtobits(-0.21613245),$shortrealtobits(0.20001395),$shortrealtobits(0.014193953),
    $shortrealtobits(-0.09715731),$shortrealtobits(-0.22626093),$shortrealtobits(0.21176445),$shortrealtobits(0.10856432),
    $shortrealtobits(0.40863353),$shortrealtobits(-0.03572945),$shortrealtobits(-0.25431183),$shortrealtobits(0.3559346),
    $shortrealtobits(0.2770792),$shortrealtobits(-0.3209043),$shortrealtobits(0.0016918648),$shortrealtobits(-0.18562572),
    $shortrealtobits(0.39714593),$shortrealtobits(-0.5636728),$shortrealtobits(-0.22676389),$shortrealtobits(0.526665),
    $shortrealtobits(0.10925218),$shortrealtobits(0.2711463),$shortrealtobits(-0.29688957),$shortrealtobits(-0.6567818),
    $shortrealtobits(0.12328347),$shortrealtobits(-0.426596),$shortrealtobits(0.4659878),$shortrealtobits(0.37539217),
    $shortrealtobits(-0.12395944),$shortrealtobits(0.35996306),$shortrealtobits(0.48443636),$shortrealtobits(0.50947547),
    $shortrealtobits(-0.28169835),$shortrealtobits(-0.32736093),$shortrealtobits(0.4576045),$shortrealtobits(0.27243197),
    $shortrealtobits(0.3658569),$shortrealtobits(-0.5254163),$shortrealtobits(0.36818987),$shortrealtobits(-0.38184917)
  },
  '{ 
    $shortrealtobits(0.18834795),$shortrealtobits(0.048145425),$shortrealtobits(-0.5607876),$shortrealtobits(0.16863126),
    $shortrealtobits(0.18892352),$shortrealtobits(-0.16903052),$shortrealtobits(-0.1850679),$shortrealtobits(0.044601902),
    $shortrealtobits(0.4626124),$shortrealtobits(0.31277362),$shortrealtobits(-0.1889117),$shortrealtobits(-0.12699938),
    $shortrealtobits(-0.15261725),$shortrealtobits(0.16448317),$shortrealtobits(0.30209482),$shortrealtobits(0.027889809),
    $shortrealtobits(0.23835334),$shortrealtobits(-0.39592728),$shortrealtobits(0.27012396),$shortrealtobits(0.44392142),
    $shortrealtobits(0.3374563),$shortrealtobits(0.3392927),$shortrealtobits(0.10233305),$shortrealtobits(-0.13167551),
    $shortrealtobits(0.13781185),$shortrealtobits(-0.5523386),$shortrealtobits(-0.35848975),$shortrealtobits(0.2529747),
    $shortrealtobits(-0.4202073),$shortrealtobits(-0.15145826),$shortrealtobits(0.49230444),$shortrealtobits(0.39031303),
    $shortrealtobits(-0.4003571),$shortrealtobits(0.4406091),$shortrealtobits(-0.13263214),$shortrealtobits(0.45968798),
    $shortrealtobits(-0.023132881),$shortrealtobits(0.3690477),$shortrealtobits(-0.4054951),$shortrealtobits(-0.04672674)
  },
  '{ 
    $shortrealtobits(-0.3013424),$shortrealtobits(0.123921014),$shortrealtobits(-0.21288301),$shortrealtobits(0.40946203),
    $shortrealtobits(-0.35644975),$shortrealtobits(-0.30458337),$shortrealtobits(0.48641518),$shortrealtobits(-0.37527254),
    $shortrealtobits(-0.040115297),$shortrealtobits(-0.17519525),$shortrealtobits(-0.4736411),$shortrealtobits(-0.3151565),
    $shortrealtobits(0.1281367),$shortrealtobits(0.07571156),$shortrealtobits(0.40711087),$shortrealtobits(-0.16408806),
    $shortrealtobits(-0.26891044),$shortrealtobits(-0.10682127),$shortrealtobits(-0.082408525),$shortrealtobits(0.22045043),
    $shortrealtobits(-0.17644002),$shortrealtobits(0.261891),$shortrealtobits(0.3143953),$shortrealtobits(-0.26342037),
    $shortrealtobits(-0.2699001),$shortrealtobits(-0.12831572),$shortrealtobits(-0.2793132),$shortrealtobits(-0.12172861),
    $shortrealtobits(0.5445982),$shortrealtobits(-0.18687035),$shortrealtobits(-0.3662606),$shortrealtobits(0.14557944),
    $shortrealtobits(0.36153704),$shortrealtobits(-0.34628958),$shortrealtobits(-0.41292298),$shortrealtobits(-0.058854517),
    $shortrealtobits(-0.3629218),$shortrealtobits(0.3071151),$shortrealtobits(0.09761916),$shortrealtobits(0.17767382)
  },
  '{ 
    $shortrealtobits(-0.12887214),$shortrealtobits(-0.26084304),$shortrealtobits(0.6695665),$shortrealtobits(-0.13954546),
    $shortrealtobits(0.43730044),$shortrealtobits(-0.5659167),$shortrealtobits(0.3385649),$shortrealtobits(0.24797846),
    $shortrealtobits(0.5555669),$shortrealtobits(-0.56024086),$shortrealtobits(0.52802145),$shortrealtobits(-0.41783533),
    $shortrealtobits(-0.28948143),$shortrealtobits(0.14119297),$shortrealtobits(0.089166574),$shortrealtobits(-0.54510194),
    $shortrealtobits(0.011694484),$shortrealtobits(-0.53716975),$shortrealtobits(0.53651565),$shortrealtobits(0.16648445),
    $shortrealtobits(0.02876113),$shortrealtobits(-0.26643872),$shortrealtobits(0.13024919),$shortrealtobits(0.7079987),
    $shortrealtobits(0.16648799),$shortrealtobits(-0.45844948),$shortrealtobits(-0.30502734),$shortrealtobits(-0.16842727),
    $shortrealtobits(0.72963077),$shortrealtobits(-0.22103353),$shortrealtobits(0.11598902),$shortrealtobits(-0.45648664),
    $shortrealtobits(0.041656584),$shortrealtobits(0.368869),$shortrealtobits(0.50761104),$shortrealtobits(-0.13356443),
    $shortrealtobits(-0.0693419),$shortrealtobits(-0.3177529),$shortrealtobits(-0.5373838),$shortrealtobits(0.5490954)
  },
  '{ 
    $shortrealtobits(0.008601378),$shortrealtobits(0.41467768),$shortrealtobits(-0.38714722),$shortrealtobits(0.32976675),
    $shortrealtobits(0.38308698),$shortrealtobits(-0.14166372),$shortrealtobits(0.34239897),$shortrealtobits(-0.089515336),
    $shortrealtobits(-0.14505455),$shortrealtobits(-0.2837298),$shortrealtobits(-0.48718217),$shortrealtobits(-0.14389166),
    $shortrealtobits(-0.30171096),$shortrealtobits(-0.24724825),$shortrealtobits(-0.15045828),$shortrealtobits(0.32971728),
    $shortrealtobits(0.2526947),$shortrealtobits(0.15553544),$shortrealtobits(-0.17721854),$shortrealtobits(0.3549754),
    $shortrealtobits(-0.00907392),$shortrealtobits(-0.1885686),$shortrealtobits(-0.07432337),$shortrealtobits(0.046408128),
    $shortrealtobits(-0.14355676),$shortrealtobits(0.43639517),$shortrealtobits(0.19867234),$shortrealtobits(-0.24290003),
    $shortrealtobits(-0.3353441),$shortrealtobits(-0.022887465),$shortrealtobits(0.10056982),$shortrealtobits(-0.29552376),
    $shortrealtobits(-0.14452904),$shortrealtobits(0.00372726),$shortrealtobits(-0.57605106),$shortrealtobits(0.003593318),
    $shortrealtobits(0.03841583),$shortrealtobits(0.3248822),$shortrealtobits(-0.03537169),$shortrealtobits(0.35257858)
  },
  '{ 
    $shortrealtobits(0.46750394),$shortrealtobits(0.20231098),$shortrealtobits(0.5038917),$shortrealtobits(0.2980287),
    $shortrealtobits(-0.29046586),$shortrealtobits(-0.10645501),$shortrealtobits(0.42859915),$shortrealtobits(0.120930456),
    $shortrealtobits(-0.08567338),$shortrealtobits(-0.19445907),$shortrealtobits(0.15881464),$shortrealtobits(0.4447534),
    $shortrealtobits(-0.23098001),$shortrealtobits(-0.34586057),$shortrealtobits(0.3527274),$shortrealtobits(0.32816646),
    $shortrealtobits(0.29186168),$shortrealtobits(-0.29679647),$shortrealtobits(0.1539707),$shortrealtobits(0.122156434),
    $shortrealtobits(0.048786525),$shortrealtobits(0.3133696),$shortrealtobits(-0.3920538),$shortrealtobits(-0.6595159),
    $shortrealtobits(-0.41268063),$shortrealtobits(0.20417576),$shortrealtobits(0.28514117),$shortrealtobits(-0.122277945),
    $shortrealtobits(0.15874447),$shortrealtobits(0.5344208),$shortrealtobits(-0.09266008),$shortrealtobits(-0.3481477),
    $shortrealtobits(-0.1695134),$shortrealtobits(-0.2534524),$shortrealtobits(0.11615478),$shortrealtobits(0.16159935),
    $shortrealtobits(0.24511723),$shortrealtobits(-0.037910435),$shortrealtobits(-0.31991225),$shortrealtobits(0.13867906)
  },
  '{ 
    $shortrealtobits(0.13155182),$shortrealtobits(0.2382443),$shortrealtobits(-0.49883682),$shortrealtobits(-0.04430887),
    $shortrealtobits(0.33066487),$shortrealtobits(-0.27564836),$shortrealtobits(-0.008740025),$shortrealtobits(0.28104514),
    $shortrealtobits(0.45177707),$shortrealtobits(-0.23850378),$shortrealtobits(-0.4481478),$shortrealtobits(0.20634782),
    $shortrealtobits(0.2930017),$shortrealtobits(0.1800656),$shortrealtobits(0.4453704),$shortrealtobits(-0.3410804),
    $shortrealtobits(-0.5172636),$shortrealtobits(0.08628713),$shortrealtobits(-0.41282007),$shortrealtobits(0.33977887),
    $shortrealtobits(-0.048518334),$shortrealtobits(-0.16198123),$shortrealtobits(0.2667012),$shortrealtobits(0.083674885),
    $shortrealtobits(-0.0030541003),$shortrealtobits(0.26411906),$shortrealtobits(-0.7496101),$shortrealtobits(0.2887101),
    $shortrealtobits(-0.5075449),$shortrealtobits(0.28055248),$shortrealtobits(-0.22446185),$shortrealtobits(0.42099822),
    $shortrealtobits(-0.2373369),$shortrealtobits(-0.021232039),$shortrealtobits(-0.49829376),$shortrealtobits(-0.4004778),
    $shortrealtobits(-0.5671661),$shortrealtobits(-0.5416571),$shortrealtobits(-0.10666899),$shortrealtobits(-0.6850164)
  },
  '{ 
    $shortrealtobits(-0.31502384),$shortrealtobits(0.3596969),$shortrealtobits(0.18136816),$shortrealtobits(0.5493342),
    $shortrealtobits(-0.36667326),$shortrealtobits(0.012407096),$shortrealtobits(0.23153253),$shortrealtobits(0.124296986),
    $shortrealtobits(-0.30231434),$shortrealtobits(-0.4049609),$shortrealtobits(0.44515774),$shortrealtobits(0.18997012),
    $shortrealtobits(0.08417451),$shortrealtobits(0.34584117),$shortrealtobits(-0.3015468),$shortrealtobits(-0.38351178),
    $shortrealtobits(0.12503713),$shortrealtobits(-0.38420793),$shortrealtobits(0.4964991),$shortrealtobits(-0.2269744),
    $shortrealtobits(0.5152238),$shortrealtobits(-0.16830826),$shortrealtobits(-0.15998723),$shortrealtobits(-0.27323252),
    $shortrealtobits(0.2508237),$shortrealtobits(0.24652225),$shortrealtobits(0.22615112),$shortrealtobits(0.23477948),
    $shortrealtobits(-0.18202685),$shortrealtobits(-0.1931531),$shortrealtobits(-0.2897782),$shortrealtobits(-0.2819795),
    $shortrealtobits(0.09315135),$shortrealtobits(-0.2502858),$shortrealtobits(-0.10046642),$shortrealtobits(0.60471296),
    $shortrealtobits(-0.39113304),$shortrealtobits(-0.065644376),$shortrealtobits(0.32999453),$shortrealtobits(0.14116026)
  },
  '{ 
    $shortrealtobits(0.61710596),$shortrealtobits(-0.32092425),$shortrealtobits(0.32451716),$shortrealtobits(-0.2042854),
    $shortrealtobits(-0.14056087),$shortrealtobits(0.0760211),$shortrealtobits(-0.53534275),$shortrealtobits(-0.06751308),
    $shortrealtobits(-0.078200996),$shortrealtobits(-0.056066502),$shortrealtobits(-0.18705487),$shortrealtobits(-0.29560643),
    $shortrealtobits(0.56478596),$shortrealtobits(-0.043562185),$shortrealtobits(0.06719454),$shortrealtobits(-0.12933095),
    $shortrealtobits(-0.22132899),$shortrealtobits(0.14653029),$shortrealtobits(0.05761323),$shortrealtobits(-0.60564226),
    $shortrealtobits(0.37257192),$shortrealtobits(0.26844606),$shortrealtobits(-0.10913576),$shortrealtobits(-0.37335378),
    $shortrealtobits(-0.3330795),$shortrealtobits(-0.4130078),$shortrealtobits(-0.010821582),$shortrealtobits(0.10691492),
    $shortrealtobits(-0.0606821),$shortrealtobits(0.17801982),$shortrealtobits(0.3025641),$shortrealtobits(0.47294345),
    $shortrealtobits(-0.46558708),$shortrealtobits(-0.30425236),$shortrealtobits(-0.75449085),$shortrealtobits(-0.059204858),
    $shortrealtobits(-0.13549697),$shortrealtobits(-0.48195925),$shortrealtobits(0.03427088),$shortrealtobits(-0.22884096)
  },
  '{ 
    $shortrealtobits(-0.24716288),$shortrealtobits(-0.006461823),$shortrealtobits(0.071802266),$shortrealtobits(0.18721563),
    $shortrealtobits(0.1513835),$shortrealtobits(-0.23725116),$shortrealtobits(-0.14933693),$shortrealtobits(0.08109586),
    $shortrealtobits(0.09930328),$shortrealtobits(-0.33007377),$shortrealtobits(0.45371148),$shortrealtobits(-0.1778533),
    $shortrealtobits(-0.3332597),$shortrealtobits(0.16677277),$shortrealtobits(-0.12506762),$shortrealtobits(0.29589424),
    $shortrealtobits(0.4458952),$shortrealtobits(0.22512443),$shortrealtobits(-0.2384671),$shortrealtobits(-0.19214551),
    $shortrealtobits(0.46270758),$shortrealtobits(0.40013677),$shortrealtobits(-0.31938794),$shortrealtobits(0.20316373),
    $shortrealtobits(-0.19688639),$shortrealtobits(0.08850655),$shortrealtobits(-0.104087986),$shortrealtobits(-0.53750324),
    $shortrealtobits(-0.17783006),$shortrealtobits(-0.09535952),$shortrealtobits(0.23423684),$shortrealtobits(-0.24475206),
    $shortrealtobits(0.08886433),$shortrealtobits(0.39555782),$shortrealtobits(0.06703721),$shortrealtobits(0.31518334),
    $shortrealtobits(0.03901229),$shortrealtobits(-0.4368169),$shortrealtobits(0.19284977),$shortrealtobits(0.058383957)
  },
  '{ 
    $shortrealtobits(-0.022070583),$shortrealtobits(-0.5526479),$shortrealtobits(0.6609293),$shortrealtobits(0.36355445),
    $shortrealtobits(-0.40992865),$shortrealtobits(-0.46491972),$shortrealtobits(-0.28429192),$shortrealtobits(-0.29278642),
    $shortrealtobits(-0.21304527),$shortrealtobits(0.12588654),$shortrealtobits(-0.34229463),$shortrealtobits(-0.0014507435),
    $shortrealtobits(-0.29045558),$shortrealtobits(-0.25428987),$shortrealtobits(0.09532856),$shortrealtobits(0.068252146),
    $shortrealtobits(-0.046394844),$shortrealtobits(-0.4561023),$shortrealtobits(0.39320898),$shortrealtobits(-0.54015404),
    $shortrealtobits(0.38906348),$shortrealtobits(0.041143406),$shortrealtobits(-0.3390535),$shortrealtobits(0.6835147),
    $shortrealtobits(-0.34022015),$shortrealtobits(-0.37564126),$shortrealtobits(0.1953739),$shortrealtobits(0.32199916),
    $shortrealtobits(0.38782188),$shortrealtobits(-0.3456122),$shortrealtobits(0.039548047),$shortrealtobits(0.4538122),
    $shortrealtobits(0.3937342),$shortrealtobits(0.033904474),$shortrealtobits(-0.536748),$shortrealtobits(-0.3442699),
    $shortrealtobits(0.19829972),$shortrealtobits(-0.44691736),$shortrealtobits(0.17009957),$shortrealtobits(-0.29609042)
  },
  '{ 
    $shortrealtobits(0.062197737),$shortrealtobits(-0.08066863),$shortrealtobits(-0.037286498),$shortrealtobits(-0.3223886),
    $shortrealtobits(0.21433382),$shortrealtobits(0.3115015),$shortrealtobits(-0.111213475),$shortrealtobits(0.22260581),
    $shortrealtobits(0.12543082),$shortrealtobits(-0.10063069),$shortrealtobits(0.06666358),$shortrealtobits(0.20371889),
    $shortrealtobits(-0.22017895),$shortrealtobits(-0.1852223),$shortrealtobits(0.27684003),$shortrealtobits(-0.036922883),
    $shortrealtobits(0.10304554),$shortrealtobits(-0.1781858),$shortrealtobits(0.09743499),$shortrealtobits(-0.15255049),
    $shortrealtobits(0.36480936),$shortrealtobits(0.45558676),$shortrealtobits(0.5001177),$shortrealtobits(-0.13704637),
    $shortrealtobits(-0.16832356),$shortrealtobits(-0.015917324),$shortrealtobits(-0.19089073),$shortrealtobits(0.019748399),
    $shortrealtobits(0.5074167),$shortrealtobits(-0.19261903),$shortrealtobits(-0.12140637),$shortrealtobits(-0.08714689),
    $shortrealtobits(-0.43684426),$shortrealtobits(-0.20417991),$shortrealtobits(0.010545772),$shortrealtobits(-0.16957045),
    $shortrealtobits(-0.4634144),$shortrealtobits(-0.633485),$shortrealtobits(-0.32882237),$shortrealtobits(0.36585373)
  },
  '{ 
    $shortrealtobits(0.24230798),$shortrealtobits(0.21859147),$shortrealtobits(-0.0022786048),$shortrealtobits(-0.04614255),
    $shortrealtobits(-0.25177753),$shortrealtobits(-0.08411275),$shortrealtobits(0.6947522),$shortrealtobits(0.42358118),
    $shortrealtobits(-0.16428412),$shortrealtobits(-0.1970231),$shortrealtobits(0.22795558),$shortrealtobits(-0.022501286),
    $shortrealtobits(-0.5042697),$shortrealtobits(0.15986843),$shortrealtobits(0.45907417),$shortrealtobits(-0.20163162),
    $shortrealtobits(0.012507349),$shortrealtobits(-0.3792546),$shortrealtobits(-0.16385663),$shortrealtobits(-0.49586508),
    $shortrealtobits(-0.3300403),$shortrealtobits(-0.40886945),$shortrealtobits(-0.1250359),$shortrealtobits(0.47042155),
    $shortrealtobits(-0.4322163),$shortrealtobits(0.31551433),$shortrealtobits(0.1964868),$shortrealtobits(0.11308127),
    $shortrealtobits(0.09023014),$shortrealtobits(0.48456037),$shortrealtobits(-0.6691253),$shortrealtobits(-0.030763231),
    $shortrealtobits(0.2005836),$shortrealtobits(-0.4035953),$shortrealtobits(-0.5840361),$shortrealtobits(0.40152687),
    $shortrealtobits(0.10580228),$shortrealtobits(-0.4347327),$shortrealtobits(-0.5739627),$shortrealtobits(0.09212967)
  },
  '{ 
    $shortrealtobits(0.3875554),$shortrealtobits(-0.044344787),$shortrealtobits(-0.19767411),$shortrealtobits(0.11191471),
    $shortrealtobits(0.28888842),$shortrealtobits(0.6367475),$shortrealtobits(-0.46705747),$shortrealtobits(-0.3490922),
    $shortrealtobits(0.14186345),$shortrealtobits(0.12131947),$shortrealtobits(-0.38523948),$shortrealtobits(-0.17567377),
    $shortrealtobits(0.34904453),$shortrealtobits(-0.39297843),$shortrealtobits(0.17238505),$shortrealtobits(-0.43874738),
    $shortrealtobits(-0.19342001),$shortrealtobits(0.37789902),$shortrealtobits(-0.04847549),$shortrealtobits(-0.3000505),
    $shortrealtobits(0.27532205),$shortrealtobits(0.09958976),$shortrealtobits(0.5455438),$shortrealtobits(0.34781176),
    $shortrealtobits(-0.03530107),$shortrealtobits(0.005462129),$shortrealtobits(0.40173537),$shortrealtobits(0.5336039),
    $shortrealtobits(-0.37862894),$shortrealtobits(0.37860546),$shortrealtobits(0.33066726),$shortrealtobits(0.42412752),
    $shortrealtobits(-0.15925045),$shortrealtobits(0.1241213),$shortrealtobits(-0.10845135),$shortrealtobits(-0.15844029),
    $shortrealtobits(0.0450602),$shortrealtobits(0.17237537),$shortrealtobits(0.04616853),$shortrealtobits(-0.31247368)
  },
  '{ 
    $shortrealtobits(-0.47936633),$shortrealtobits(0.060117543),$shortrealtobits(-0.062148772),$shortrealtobits(-0.26793745),
    $shortrealtobits(-0.49341065),$shortrealtobits(-0.4588345),$shortrealtobits(-0.18353255),$shortrealtobits(-0.3447495),
    $shortrealtobits(0.02348414),$shortrealtobits(-0.7102928),$shortrealtobits(0.31979248),$shortrealtobits(-0.10536521),
    $shortrealtobits(-0.17182027),$shortrealtobits(-0.30473378),$shortrealtobits(0.021064574),$shortrealtobits(-0.32371047),
    $shortrealtobits(-0.03219028),$shortrealtobits(0.30231428),$shortrealtobits(0.4389021),$shortrealtobits(0.34703785),
    $shortrealtobits(0.3772842),$shortrealtobits(0.27504915),$shortrealtobits(0.27567348),$shortrealtobits(-0.3281041),
    $shortrealtobits(-0.007547174),$shortrealtobits(0.03454182),$shortrealtobits(0.22622181),$shortrealtobits(0.46550983),
    $shortrealtobits(0.060201056),$shortrealtobits(0.39042696),$shortrealtobits(0.6406243),$shortrealtobits(0.17523539),
    $shortrealtobits(-0.3720006),$shortrealtobits(-0.32774544),$shortrealtobits(0.07093173),$shortrealtobits(-0.20455031),
    $shortrealtobits(-0.5949119),$shortrealtobits(0.22594975),$shortrealtobits(0.06765888),$shortrealtobits(-0.25673643)
  },
  '{ 
    $shortrealtobits(-0.25855803),$shortrealtobits(0.048261702),$shortrealtobits(-0.37120345),$shortrealtobits(0.1516445),
    $shortrealtobits(-0.6562714),$shortrealtobits(-0.7137253),$shortrealtobits(0.26928982),$shortrealtobits(-0.4272919),
    $shortrealtobits(-0.585662),$shortrealtobits(-0.21888772),$shortrealtobits(-0.1370984),$shortrealtobits(-0.10724953),
    $shortrealtobits(-0.054714467),$shortrealtobits(0.5903472),$shortrealtobits(0.04164072),$shortrealtobits(-0.15217459),
    $shortrealtobits(0.3891272),$shortrealtobits(-0.27601954),$shortrealtobits(0.022649778),$shortrealtobits(-0.3121524),
    $shortrealtobits(-0.10199726),$shortrealtobits(0.4123153),$shortrealtobits(-0.13332357),$shortrealtobits(0.47253838),
    $shortrealtobits(0.16375698),$shortrealtobits(-0.4104111),$shortrealtobits(-0.46332803),$shortrealtobits(-0.20098104),
    $shortrealtobits(0.25428364),$shortrealtobits(0.37802127),$shortrealtobits(-0.3538325),$shortrealtobits(0.090763986),
    $shortrealtobits(0.07850684),$shortrealtobits(-0.102113724),$shortrealtobits(0.27553043),$shortrealtobits(0.045995314),
    $shortrealtobits(0.35208422),$shortrealtobits(-0.31511113),$shortrealtobits(0.44448695),$shortrealtobits(-0.41566512)
  },
  '{ 
    $shortrealtobits(-0.09128631),$shortrealtobits(-0.26657233),$shortrealtobits(0.38950288),$shortrealtobits(-0.028712573),
    $shortrealtobits(0.08992213),$shortrealtobits(-0.46933764),$shortrealtobits(-0.23614214),$shortrealtobits(0.3226318),
    $shortrealtobits(-0.10399784),$shortrealtobits(0.29240185),$shortrealtobits(0.5919349),$shortrealtobits(0.42732623),
    $shortrealtobits(-0.3624164),$shortrealtobits(-0.12308498),$shortrealtobits(-0.44457036),$shortrealtobits(0.37856314),
    $shortrealtobits(-0.19827098),$shortrealtobits(0.017271515),$shortrealtobits(0.13028757),$shortrealtobits(-0.36618164),
    $shortrealtobits(-0.39966875),$shortrealtobits(0.22228956),$shortrealtobits(-0.21488222),$shortrealtobits(0.23386759),
    $shortrealtobits(-0.40143117),$shortrealtobits(0.086719945),$shortrealtobits(-0.41953242),$shortrealtobits(-0.10062717),
    $shortrealtobits(-0.07591705),$shortrealtobits(-0.30223462),$shortrealtobits(-0.009523059),$shortrealtobits(-0.44885254),
    $shortrealtobits(0.12018305),$shortrealtobits(0.25384846),$shortrealtobits(-0.4705305),$shortrealtobits(-0.5129938),
    $shortrealtobits(-0.08488335),$shortrealtobits(-0.33417973),$shortrealtobits(0.043593667),$shortrealtobits(-0.39038482)
  },
  '{ 
    $shortrealtobits(0.35228977),$shortrealtobits(-0.024619883),$shortrealtobits(0.1578588),$shortrealtobits(-0.11478718),
    $shortrealtobits(-0.12284468),$shortrealtobits(0.15569027),$shortrealtobits(0.023563432),$shortrealtobits(-0.24659267),
    $shortrealtobits(0.37286508),$shortrealtobits(0.025921347),$shortrealtobits(0.2872955),$shortrealtobits(0.37136188),
    $shortrealtobits(-0.4225257),$shortrealtobits(-0.2034195),$shortrealtobits(-0.34613863),$shortrealtobits(-0.28452736),
    $shortrealtobits(0.769043),$shortrealtobits(-0.22985885),$shortrealtobits(-0.017530201),$shortrealtobits(-0.18670522),
    $shortrealtobits(-0.039962325),$shortrealtobits(-0.2984973),$shortrealtobits(-0.105492234),$shortrealtobits(-0.28299877),
    $shortrealtobits(-0.2363268),$shortrealtobits(0.2150083),$shortrealtobits(-0.21875653),$shortrealtobits(-0.87831837),
    $shortrealtobits(-0.32586145),$shortrealtobits(0.31295085),$shortrealtobits(-0.9630084),$shortrealtobits(-0.026971726),
    $shortrealtobits(-0.40192506),$shortrealtobits(-0.19278762),$shortrealtobits(0.13623972),$shortrealtobits(0.16542535),
    $shortrealtobits(0.024087034),$shortrealtobits(0.058380492),$shortrealtobits(-0.29023224),$shortrealtobits(0.14438604)
  },
  '{ 
    $shortrealtobits(-0.044594765),$shortrealtobits(-0.11703816),$shortrealtobits(0.5038497),$shortrealtobits(-0.3416401),
    $shortrealtobits(-0.65437424),$shortrealtobits(-0.44404647),$shortrealtobits(0.21142471),$shortrealtobits(0.013325923),
    $shortrealtobits(0.19515698),$shortrealtobits(0.14420418),$shortrealtobits(-0.13675962),$shortrealtobits(-0.34791112),
    $shortrealtobits(-0.42948186),$shortrealtobits(-0.044209916),$shortrealtobits(-0.4143781),$shortrealtobits(0.11053111),
    $shortrealtobits(-0.16039552),$shortrealtobits(-0.3973279),$shortrealtobits(0.27889594),$shortrealtobits(-0.30919233),
    $shortrealtobits(-0.31563434),$shortrealtobits(0.41558668),$shortrealtobits(-0.12823686),$shortrealtobits(-0.10995439),
    $shortrealtobits(-0.5268131),$shortrealtobits(-0.113457),$shortrealtobits(-0.2533313),$shortrealtobits(-0.49784777),
    $shortrealtobits(-0.073486544),$shortrealtobits(0.006993058),$shortrealtobits(0.15584698),$shortrealtobits(0.22353166),
    $shortrealtobits(0.3939995),$shortrealtobits(-0.15587151),$shortrealtobits(0.17189872),$shortrealtobits(-0.32287544),
    $shortrealtobits(-0.20981146),$shortrealtobits(-0.30048203),$shortrealtobits(-0.32107866),$shortrealtobits(-0.21535772)
  },
  '{ 
    $shortrealtobits(-0.49149922),$shortrealtobits(-0.31346974),$shortrealtobits(0.15210983),$shortrealtobits(0.34554106),
    $shortrealtobits(-0.18316585),$shortrealtobits(-0.43158615),$shortrealtobits(0.09165978),$shortrealtobits(0.30436045),
    $shortrealtobits(-0.41404507),$shortrealtobits(-0.121041715),$shortrealtobits(0.29622382),$shortrealtobits(-0.29498282),
    $shortrealtobits(-0.37830332),$shortrealtobits(0.5550934),$shortrealtobits(-0.039658513),$shortrealtobits(-0.070796564),
    $shortrealtobits(0.5614065),$shortrealtobits(-0.3648446),$shortrealtobits(-0.062883414),$shortrealtobits(-0.3133227),
    $shortrealtobits(0.30331177),$shortrealtobits(-0.27915812),$shortrealtobits(-0.05741999),$shortrealtobits(0.11794625),
    $shortrealtobits(0.3704765),$shortrealtobits(0.10342637),$shortrealtobits(0.11853399),$shortrealtobits(0.40283912),
    $shortrealtobits(-0.24324507),$shortrealtobits(-0.16693974),$shortrealtobits(-0.32849672),$shortrealtobits(-0.027752804),
    $shortrealtobits(0.17361341),$shortrealtobits(-0.39704195),$shortrealtobits(0.23901455),$shortrealtobits(-0.16846277),
    $shortrealtobits(0.5266464),$shortrealtobits(-0.121081375),$shortrealtobits(-0.20892705),$shortrealtobits(-0.098624825)
  },
  '{ 
    $shortrealtobits(0.22704835),$shortrealtobits(-0.44491753),$shortrealtobits(0.8128013),$shortrealtobits(0.49257722),
    $shortrealtobits(-0.022706004),$shortrealtobits(-0.36971548),$shortrealtobits(0.32686204),$shortrealtobits(0.06410507),
    $shortrealtobits(-0.34425238),$shortrealtobits(0.47516346),$shortrealtobits(0.34729394),$shortrealtobits(-0.29141912),
    $shortrealtobits(0.12690865),$shortrealtobits(-0.1546628),$shortrealtobits(0.06728576),$shortrealtobits(-0.13909997),
    $shortrealtobits(-0.281431),$shortrealtobits(0.24412489),$shortrealtobits(0.2883115),$shortrealtobits(-0.28107557),
    $shortrealtobits(0.39464492),$shortrealtobits(-0.41282043),$shortrealtobits(-0.28547114),$shortrealtobits(0.37875354),
    $shortrealtobits(0.27009606),$shortrealtobits(-0.08827446),$shortrealtobits(-0.27287033),$shortrealtobits(-0.72494644),
    $shortrealtobits(-0.54001117),$shortrealtobits(0.14942178),$shortrealtobits(0.022237659),$shortrealtobits(-0.4451745),
    $shortrealtobits(0.21948232),$shortrealtobits(0.33659592),$shortrealtobits(-0.1623364),$shortrealtobits(-0.08701209),
    $shortrealtobits(-0.43912244),$shortrealtobits(-0.33601254),$shortrealtobits(-0.427094),$shortrealtobits(-0.31990007)
  },
  '{ 
    $shortrealtobits(0.5445667),$shortrealtobits(-0.12711684),$shortrealtobits(0.40735486),$shortrealtobits(-0.27956417),
    $shortrealtobits(-0.09775135),$shortrealtobits(-0.17655273),$shortrealtobits(0.10259035),$shortrealtobits(0.23491882),
    $shortrealtobits(-0.6791216),$shortrealtobits(0.78641284),$shortrealtobits(0.33858758),$shortrealtobits(0.48976868),
    $shortrealtobits(-0.48245364),$shortrealtobits(-0.056096613),$shortrealtobits(-0.015717143),$shortrealtobits(0.44485423),
    $shortrealtobits(0.05817248),$shortrealtobits(-0.16373357),$shortrealtobits(0.13167138),$shortrealtobits(-0.33188123),
    $shortrealtobits(0.4273957),$shortrealtobits(0.30858088),$shortrealtobits(-0.3208396),$shortrealtobits(0.7005892),
    $shortrealtobits(0.33862904),$shortrealtobits(0.28182742),$shortrealtobits(0.30795327),$shortrealtobits(0.43567336),
    $shortrealtobits(-0.3974354),$shortrealtobits(-0.2584003),$shortrealtobits(0.032559354),$shortrealtobits(-0.06348215),
    $shortrealtobits(0.32872924),$shortrealtobits(-0.07222894),$shortrealtobits(0.5030089),$shortrealtobits(-0.15250282),
    $shortrealtobits(0.5679436),$shortrealtobits(0.18298988),$shortrealtobits(-0.6990384),$shortrealtobits(-0.42974707)
  },
  '{ 
    $shortrealtobits(0.5571906),$shortrealtobits(-0.03258611),$shortrealtobits(0.36959764),$shortrealtobits(0.3493097),
    $shortrealtobits(-0.38977802),$shortrealtobits(0.2238102),$shortrealtobits(0.1278121),$shortrealtobits(0.14971523),
    $shortrealtobits(0.034696043),$shortrealtobits(-0.35132626),$shortrealtobits(-0.33335483),$shortrealtobits(-0.39236608),
    $shortrealtobits(0.25818163),$shortrealtobits(0.36405742),$shortrealtobits(0.26089564),$shortrealtobits(0.2616201),
    $shortrealtobits(-0.5562446),$shortrealtobits(-0.011215636),$shortrealtobits(0.35617712),$shortrealtobits(0.08709058),
    $shortrealtobits(0.24440347),$shortrealtobits(-0.029730532),$shortrealtobits(-0.15590844),$shortrealtobits(0.42303666),
    $shortrealtobits(-0.07196841),$shortrealtobits(-0.008128353),$shortrealtobits(-0.7718027),$shortrealtobits(0.051972367),
    $shortrealtobits(-0.04930397),$shortrealtobits(0.46990106),$shortrealtobits(-0.05220313),$shortrealtobits(-0.20446175),
    $shortrealtobits(-0.49944136),$shortrealtobits(0.3272594),$shortrealtobits(-0.5026745),$shortrealtobits(-0.33509523),
    $shortrealtobits(-0.15497686),$shortrealtobits(-0.09329873),$shortrealtobits(0.0054774224),$shortrealtobits(-0.7026961)
  },
  '{ 
    $shortrealtobits(0.2756096),$shortrealtobits(0.1700448),$shortrealtobits(0.29026124),$shortrealtobits(-0.4236831),
    $shortrealtobits(0.12937029),$shortrealtobits(-0.03735541),$shortrealtobits(-0.08915504),$shortrealtobits(0.47072273),
    $shortrealtobits(0.172436),$shortrealtobits(0.42853686),$shortrealtobits(0.058185678),$shortrealtobits(0.47163242),
    $shortrealtobits(0.3039216),$shortrealtobits(0.12715058),$shortrealtobits(-0.08191338),$shortrealtobits(-0.35300186),
    $shortrealtobits(-0.24027379),$shortrealtobits(-0.32607663),$shortrealtobits(-0.38947412),$shortrealtobits(-0.4300698),
    $shortrealtobits(0.43113792),$shortrealtobits(0.25257802),$shortrealtobits(0.16914079),$shortrealtobits(0.50174385),
    $shortrealtobits(-0.2086651),$shortrealtobits(-0.3184383),$shortrealtobits(-0.21827547),$shortrealtobits(0.07044553),
    $shortrealtobits(0.3484614),$shortrealtobits(0.3853309),$shortrealtobits(-0.011660298),$shortrealtobits(-0.151368),
    $shortrealtobits(0.061827242),$shortrealtobits(0.20958722),$shortrealtobits(-0.31778398),$shortrealtobits(-0.41479942),
    $shortrealtobits(-0.08223102),$shortrealtobits(-0.2631226),$shortrealtobits(-0.1827484),$shortrealtobits(0.029364802)
  },
  '{ 
    $shortrealtobits(0.13729389),$shortrealtobits(0.3498742),$shortrealtobits(0.078668654),$shortrealtobits(-0.5363253),
    $shortrealtobits(-0.19626276),$shortrealtobits(0.24562381),$shortrealtobits(-0.30833077),$shortrealtobits(0.18297839),
    $shortrealtobits(0.061841525),$shortrealtobits(-0.07576932),$shortrealtobits(0.2623622),$shortrealtobits(-0.11655393),
    $shortrealtobits(0.15074687),$shortrealtobits(0.13102435),$shortrealtobits(-0.49471962),$shortrealtobits(-0.27428082),
    $shortrealtobits(0.14905795),$shortrealtobits(0.051212166),$shortrealtobits(0.3093746),$shortrealtobits(0.100204736),
    $shortrealtobits(-0.043999743),$shortrealtobits(0.23629251),$shortrealtobits(-0.08208317),$shortrealtobits(-0.30433366),
    $shortrealtobits(-0.24004419),$shortrealtobits(0.15754114),$shortrealtobits(-0.18762664),$shortrealtobits(0.54888856),
    $shortrealtobits(0.04567012),$shortrealtobits(-0.21603344),$shortrealtobits(-0.6494505),$shortrealtobits(0.42968056),
    $shortrealtobits(-0.070877284),$shortrealtobits(-0.43562618),$shortrealtobits(0.3958578),$shortrealtobits(-0.5069829),
    $shortrealtobits(0.3346145),$shortrealtobits(-0.030636473),$shortrealtobits(0.15561755),$shortrealtobits(-0.4323146)
  },
  '{ 
    $shortrealtobits(0.18016389),$shortrealtobits(-0.46594837),$shortrealtobits(-0.09318007),$shortrealtobits(0.0058390894),
    $shortrealtobits(0.31581575),$shortrealtobits(0.4215426),$shortrealtobits(0.18929419),$shortrealtobits(-0.3376778),
    $shortrealtobits(0.15582663),$shortrealtobits(0.32626957),$shortrealtobits(-0.26871464),$shortrealtobits(0.012258524),
    $shortrealtobits(-0.043543562),$shortrealtobits(0.2940275),$shortrealtobits(0.20144148),$shortrealtobits(0.07553021),
    $shortrealtobits(-0.4242509),$shortrealtobits(-0.1164276),$shortrealtobits(-0.24700318),$shortrealtobits(0.072904274),
    $shortrealtobits(0.20129052),$shortrealtobits(0.49152938),$shortrealtobits(0.12830873),$shortrealtobits(0.25939357),
    $shortrealtobits(0.35727245),$shortrealtobits(0.20452441),$shortrealtobits(-0.1217134),$shortrealtobits(0.049476206),
    $shortrealtobits(0.6131289),$shortrealtobits(0.013846406),$shortrealtobits(0.2307264),$shortrealtobits(0.4722143),
    $shortrealtobits(-0.3370059),$shortrealtobits(0.39177462),$shortrealtobits(-0.8712984),$shortrealtobits(-0.15915486),
    $shortrealtobits(0.21599543),$shortrealtobits(-0.1931951),$shortrealtobits(0.46048254),$shortrealtobits(-0.20963101)
  },
  '{ 
    $shortrealtobits(0.46377522),$shortrealtobits(-0.018912818),$shortrealtobits(0.105668485),$shortrealtobits(-0.0406002),
    $shortrealtobits(0.12125695),$shortrealtobits(0.12811631),$shortrealtobits(0.51306283),$shortrealtobits(-0.38390997),
    $shortrealtobits(0.14005674),$shortrealtobits(0.4853098),$shortrealtobits(0.5247326),$shortrealtobits(-0.08485374),
    $shortrealtobits(-0.037317216),$shortrealtobits(0.42226878),$shortrealtobits(-0.33909804),$shortrealtobits(0.05667284),
    $shortrealtobits(-0.11689721),$shortrealtobits(-0.28583622),$shortrealtobits(0.4599401),$shortrealtobits(-0.23796248),
    $shortrealtobits(0.42742556),$shortrealtobits(-0.066983745),$shortrealtobits(0.3095217),$shortrealtobits(-0.38170815),
    $shortrealtobits(-0.43174967),$shortrealtobits(-0.22577488),$shortrealtobits(-0.39519206),$shortrealtobits(0.15269724),
    $shortrealtobits(-0.20715114),$shortrealtobits(0.38378873),$shortrealtobits(-0.015808536),$shortrealtobits(-0.047429923),
    $shortrealtobits(0.22777005),$shortrealtobits(-0.14161146),$shortrealtobits(-0.09501042),$shortrealtobits(0.065989636),
    $shortrealtobits(-0.10368182),$shortrealtobits(-0.2751146),$shortrealtobits(-0.49015474),$shortrealtobits(0.10879558)
  },
  '{ 
    $shortrealtobits(-0.14652954),$shortrealtobits(-0.007266439),$shortrealtobits(-0.15900116),$shortrealtobits(0.54582584),
    $shortrealtobits(-0.20498337),$shortrealtobits(0.46108606),$shortrealtobits(-0.057960346),$shortrealtobits(-0.08368445),
    $shortrealtobits(-0.21290208),$shortrealtobits(0.4738483),$shortrealtobits(0.49858657),$shortrealtobits(-0.09359919),
    $shortrealtobits(0.1603282),$shortrealtobits(-0.06946713),$shortrealtobits(-0.29415667),$shortrealtobits(-0.17517579),
    $shortrealtobits(-0.30692086),$shortrealtobits(-0.097036175),$shortrealtobits(-0.0012150595),$shortrealtobits(-0.25720322),
    $shortrealtobits(0.06359598),$shortrealtobits(0.29901403),$shortrealtobits(-0.23720282),$shortrealtobits(0.53462785),
    $shortrealtobits(0.5386858),$shortrealtobits(0.22504598),$shortrealtobits(-0.5004932),$shortrealtobits(0.056442514),
    $shortrealtobits(0.16587798),$shortrealtobits(-0.06903721),$shortrealtobits(0.65500236),$shortrealtobits(0.26634616),
    $shortrealtobits(-0.49244112),$shortrealtobits(0.111918114),$shortrealtobits(0.017682374),$shortrealtobits(0.1302335),
    $shortrealtobits(0.04008827),$shortrealtobits(0.25724855),$shortrealtobits(0.0714029),$shortrealtobits(0.33872962)
  },
  '{ 
    $shortrealtobits(-0.33546627),$shortrealtobits(-0.188096),$shortrealtobits(-0.004801139),$shortrealtobits(-0.098383024),
    $shortrealtobits(0.28295213),$shortrealtobits(-0.08091173),$shortrealtobits(-0.7894826),$shortrealtobits(0.33206302),
    $shortrealtobits(-0.050734095),$shortrealtobits(0.18351783),$shortrealtobits(0.18389934),$shortrealtobits(-0.17628445),
    $shortrealtobits(0.15996592),$shortrealtobits(-0.4793298),$shortrealtobits(-0.34351325),$shortrealtobits(-0.39596325),
    $shortrealtobits(-0.27756518),$shortrealtobits(-0.2272024),$shortrealtobits(-0.12611122),$shortrealtobits(0.05448954),
    $shortrealtobits(-0.0864904),$shortrealtobits(0.019309357),$shortrealtobits(0.07664264),$shortrealtobits(0.20792106),
    $shortrealtobits(-0.26822522),$shortrealtobits(0.018640056),$shortrealtobits(0.14819378),$shortrealtobits(0.22687103),
    $shortrealtobits(0.3204357),$shortrealtobits(-0.22793445),$shortrealtobits(0.4722776),$shortrealtobits(-0.07558816),
    $shortrealtobits(0.3958265),$shortrealtobits(0.46266967),$shortrealtobits(-0.6351403),$shortrealtobits(0.43223932),
    $shortrealtobits(-0.6021805),$shortrealtobits(0.3405321),$shortrealtobits(0.02482756),$shortrealtobits(-0.19725734)
  },
  '{ 
    $shortrealtobits(-0.17912154),$shortrealtobits(-0.3414342),$shortrealtobits(0.40597922),$shortrealtobits(0.40517488),
    $shortrealtobits(-0.03527555),$shortrealtobits(-0.0021558872),$shortrealtobits(-0.6452283),$shortrealtobits(0.050333116),
    $shortrealtobits(-0.48495337),$shortrealtobits(-0.2966545),$shortrealtobits(-0.34513584),$shortrealtobits(0.106715634),
    $shortrealtobits(0.035289604),$shortrealtobits(0.017084735),$shortrealtobits(-0.14113694),$shortrealtobits(-0.5095245),
    $shortrealtobits(-0.11785698),$shortrealtobits(-0.5133703),$shortrealtobits(0.40646482),$shortrealtobits(0.10366761),
    $shortrealtobits(-0.2624869),$shortrealtobits(-0.094548784),$shortrealtobits(0.33366373),$shortrealtobits(0.59434694),
    $shortrealtobits(-0.23606388),$shortrealtobits(-0.09054527),$shortrealtobits(0.40501082),$shortrealtobits(0.457019),
    $shortrealtobits(-0.66499305),$shortrealtobits(-0.048509087),$shortrealtobits(0.77191174),$shortrealtobits(0.28777033),
    $shortrealtobits(-0.090836555),$shortrealtobits(0.21222149),$shortrealtobits(0.4294015),$shortrealtobits(-0.31287056),
    $shortrealtobits(0.47402936),$shortrealtobits(-0.22286017),$shortrealtobits(-0.17386208),$shortrealtobits(-0.006092323)
  },
  '{ 
    $shortrealtobits(-0.19382754),$shortrealtobits(0.3620087),$shortrealtobits(-0.6110025),$shortrealtobits(0.443968),
    $shortrealtobits(0.056021713),$shortrealtobits(0.6873028),$shortrealtobits(0.43094608),$shortrealtobits(0.16860008),
    $shortrealtobits(-0.11770552),$shortrealtobits(0.415552),$shortrealtobits(-0.06562017),$shortrealtobits(-0.27690598),
    $shortrealtobits(0.26098946),$shortrealtobits(-0.024129393),$shortrealtobits(0.6005215),$shortrealtobits(0.12452559),
    $shortrealtobits(-0.4532074),$shortrealtobits(0.26993805),$shortrealtobits(-0.16180024),$shortrealtobits(0.55506235),
    $shortrealtobits(0.23108195),$shortrealtobits(0.3980448),$shortrealtobits(0.3614711),$shortrealtobits(0.18111488),
    $shortrealtobits(-0.14847803),$shortrealtobits(-0.2089521),$shortrealtobits(-0.049941868),$shortrealtobits(0.6132599),
    $shortrealtobits(0.0904857),$shortrealtobits(-0.0796373),$shortrealtobits(0.021910476),$shortrealtobits(0.5112441),
    $shortrealtobits(0.37789056),$shortrealtobits(0.31799006),$shortrealtobits(-0.4617557),$shortrealtobits(0.118210025),
    $shortrealtobits(0.6173336),$shortrealtobits(-0.67985916),$shortrealtobits(-0.15453526),$shortrealtobits(0.22522676)
  },
  '{ 
    $shortrealtobits(-0.27286103),$shortrealtobits(0.38698804),$shortrealtobits(0.7050422),$shortrealtobits(-0.12505749),
    $shortrealtobits(-0.4716394),$shortrealtobits(0.045822542),$shortrealtobits(-0.44609874),$shortrealtobits(-0.1516447),
    $shortrealtobits(0.48957145),$shortrealtobits(-0.60548705),$shortrealtobits(0.16398653),$shortrealtobits(-0.3596885),
    $shortrealtobits(-0.0928979),$shortrealtobits(0.30462065),$shortrealtobits(-0.24430162),$shortrealtobits(-0.34395108),
    $shortrealtobits(0.20514035),$shortrealtobits(-0.04982454),$shortrealtobits(-0.44275558),$shortrealtobits(0.079732634),
    $shortrealtobits(-0.18660969),$shortrealtobits(-0.26243848),$shortrealtobits(-0.36680087),$shortrealtobits(0.034959532),
    $shortrealtobits(-0.47154915),$shortrealtobits(-0.30019715),$shortrealtobits(-0.130648),$shortrealtobits(-0.07991244),
    $shortrealtobits(-0.19272101),$shortrealtobits(0.67832714),$shortrealtobits(-0.09516192),$shortrealtobits(-0.47917068),
    $shortrealtobits(0.091877736),$shortrealtobits(0.1109611),$shortrealtobits(0.54856265),$shortrealtobits(-0.3489213),
    $shortrealtobits(-0.16192335),$shortrealtobits(0.012366924),$shortrealtobits(0.015401364),$shortrealtobits(-0.1965331)
  },
  '{ 
    $shortrealtobits(0.09106364),$shortrealtobits(-0.10650167),$shortrealtobits(0.3015615),$shortrealtobits(-0.3159559),
    $shortrealtobits(-0.069126524),$shortrealtobits(0.15976198),$shortrealtobits(-0.381118),$shortrealtobits(-0.12543035),
    $shortrealtobits(-0.14090511),$shortrealtobits(0.23594046),$shortrealtobits(0.2776267),$shortrealtobits(-0.0147768445),
    $shortrealtobits(0.25790703),$shortrealtobits(-0.3552054),$shortrealtobits(-0.039702304),$shortrealtobits(-0.26028103),
    $shortrealtobits(-0.39567634),$shortrealtobits(0.15885335),$shortrealtobits(0.01349335),$shortrealtobits(-0.034423634),
    $shortrealtobits(-0.08464884),$shortrealtobits(-0.34826642),$shortrealtobits(0.15319479),$shortrealtobits(-0.21825607),
    $shortrealtobits(0.3098702),$shortrealtobits(-0.407193),$shortrealtobits(-0.09622988),$shortrealtobits(0.31459555),
    $shortrealtobits(-0.5085116),$shortrealtobits(0.6358216),$shortrealtobits(0.22881663),$shortrealtobits(-0.3262676),
    $shortrealtobits(0.00802141),$shortrealtobits(0.24049035),$shortrealtobits(0.2995618),$shortrealtobits(-0.1869221),
    $shortrealtobits(0.62831455),$shortrealtobits(0.7034608),$shortrealtobits(-0.38395497),$shortrealtobits(0.64706147)
  },
  '{ 
    $shortrealtobits(0.36742425),$shortrealtobits(-0.14983332),$shortrealtobits(0.56503224),$shortrealtobits(0.3013965),
    $shortrealtobits(0.120631166),$shortrealtobits(0.093140766),$shortrealtobits(-0.254018),$shortrealtobits(0.5000985),
    $shortrealtobits(0.025628902),$shortrealtobits(0.11344145),$shortrealtobits(0.10834068),$shortrealtobits(0.5883652),
    $shortrealtobits(-0.13547875),$shortrealtobits(0.49601117),$shortrealtobits(0.22622779),$shortrealtobits(0.2966918),
    $shortrealtobits(0.37396523),$shortrealtobits(-0.3774757),$shortrealtobits(0.29955435),$shortrealtobits(0.16358727),
    $shortrealtobits(0.057191983),$shortrealtobits(-0.3327944),$shortrealtobits(0.16135831),$shortrealtobits(0.0570774),
    $shortrealtobits(0.34229815),$shortrealtobits(0.013025384),$shortrealtobits(0.40154392),$shortrealtobits(-0.06905044),
    $shortrealtobits(0.030325234),$shortrealtobits(-0.36621904),$shortrealtobits(-0.084896736),$shortrealtobits(-0.47487503),
    $shortrealtobits(-0.3059938),$shortrealtobits(-0.011626218),$shortrealtobits(0.36610022),$shortrealtobits(-0.5144629),
    $shortrealtobits(-0.14905375),$shortrealtobits(-0.28013143),$shortrealtobits(-0.027063968),$shortrealtobits(-0.46571898)
  },
  '{ 
    $shortrealtobits(-0.39828783),$shortrealtobits(0.043900643),$shortrealtobits(-0.5885966),$shortrealtobits(-0.29583618),
    $shortrealtobits(0.49107057),$shortrealtobits(0.41332275),$shortrealtobits(0.519792),$shortrealtobits(0.22824554),
    $shortrealtobits(0.27293268),$shortrealtobits(0.06717153),$shortrealtobits(-0.27146682),$shortrealtobits(-0.17494157),
    $shortrealtobits(-0.014616594),$shortrealtobits(-0.36717924),$shortrealtobits(-0.016060479),$shortrealtobits(-0.30462208),
    $shortrealtobits(0.09308992),$shortrealtobits(0.090900056),$shortrealtobits(0.07870368),$shortrealtobits(-0.05768064),
    $shortrealtobits(0.23459893),$shortrealtobits(-0.25713423),$shortrealtobits(-0.3672294),$shortrealtobits(-0.20348498),
    $shortrealtobits(0.23418666),$shortrealtobits(-0.33735177),$shortrealtobits(0.04598545),$shortrealtobits(-0.28193015),
    $shortrealtobits(0.039691657),$shortrealtobits(0.23846345),$shortrealtobits(-0.15968733),$shortrealtobits(0.34522218),
    $shortrealtobits(-0.23622242),$shortrealtobits(0.28132787),$shortrealtobits(-0.3509961),$shortrealtobits(0.16256338),
    $shortrealtobits(-0.11956838),$shortrealtobits(0.33543178),$shortrealtobits(0.7598711),$shortrealtobits(-0.12739614)
  },
  '{ 
    $shortrealtobits(-0.5925221),$shortrealtobits(0.013152432),$shortrealtobits(0.31499726),$shortrealtobits(-0.428975),
    $shortrealtobits(0.014330272),$shortrealtobits(-0.18249285),$shortrealtobits(-0.3582768),$shortrealtobits(0.53405),
    $shortrealtobits(-0.16122136),$shortrealtobits(0.43097687),$shortrealtobits(0.51787853),$shortrealtobits(0.42795128),
    $shortrealtobits(0.33632138),$shortrealtobits(-0.23078296),$shortrealtobits(-0.21458125),$shortrealtobits(0.18527362),
    $shortrealtobits(0.3158108),$shortrealtobits(0.0916335),$shortrealtobits(-0.3235685),$shortrealtobits(-0.9128643),
    $shortrealtobits(0.18533102),$shortrealtobits(0.18929385),$shortrealtobits(0.42411175),$shortrealtobits(0.66266775),
    $shortrealtobits(0.42186794),$shortrealtobits(0.19198886),$shortrealtobits(0.13676174),$shortrealtobits(-0.10395715),
    $shortrealtobits(-0.25507194),$shortrealtobits(0.012034251),$shortrealtobits(0.2647647),$shortrealtobits(0.21414147),
    $shortrealtobits(-0.3978085),$shortrealtobits(-0.39264196),$shortrealtobits(-0.42399958),$shortrealtobits(0.1405739),
    $shortrealtobits(-0.12199655),$shortrealtobits(-0.23817821),$shortrealtobits(-0.5682998),$shortrealtobits(0.30095005)
  },
  '{ 
    $shortrealtobits(0.6051671),$shortrealtobits(0.061375257),$shortrealtobits(-0.014777524),$shortrealtobits(0.3711529),
    $shortrealtobits(-0.65150505),$shortrealtobits(0.3473093),$shortrealtobits(-0.44839174),$shortrealtobits(-0.44195586),
    $shortrealtobits(-0.613537),$shortrealtobits(0.35285547),$shortrealtobits(-0.41538545),$shortrealtobits(-0.3789332),
    $shortrealtobits(0.45634872),$shortrealtobits(0.002857248),$shortrealtobits(-0.07591157),$shortrealtobits(0.3792604),
    $shortrealtobits(-0.25965214),$shortrealtobits(0.497154),$shortrealtobits(0.055349715),$shortrealtobits(0.4421081),
    $shortrealtobits(-0.19344501),$shortrealtobits(-0.04389182),$shortrealtobits(-0.1349812),$shortrealtobits(0.5012922),
    $shortrealtobits(-0.53919905),$shortrealtobits(0.46749023),$shortrealtobits(-0.012095028),$shortrealtobits(0.43372148),
    $shortrealtobits(-0.27220127),$shortrealtobits(0.3937549),$shortrealtobits(0.074489176),$shortrealtobits(0.03684331),
    $shortrealtobits(-0.23751566),$shortrealtobits(-0.097015984),$shortrealtobits(0.23439474),$shortrealtobits(0.09620926),
    $shortrealtobits(0.31423163),$shortrealtobits(0.04812298),$shortrealtobits(-0.42395353),$shortrealtobits(-0.5829853)
  },
  '{ 
    $shortrealtobits(-0.043474928),$shortrealtobits(0.119931325),$shortrealtobits(-0.1350249),$shortrealtobits(-0.32002363),
    $shortrealtobits(-0.32578805),$shortrealtobits(-0.30467165),$shortrealtobits(0.120453715),$shortrealtobits(-0.2809885),
    $shortrealtobits(-0.29791975),$shortrealtobits(-0.18988757),$shortrealtobits(0.005407705),$shortrealtobits(0.41185942),
    $shortrealtobits(0.045321018),$shortrealtobits(-0.1406978),$shortrealtobits(-0.10414728),$shortrealtobits(-0.3169139),
    $shortrealtobits(-0.19543087),$shortrealtobits(-0.31000492),$shortrealtobits(-0.27487212),$shortrealtobits(-0.35040873),
    $shortrealtobits(-0.5989894),$shortrealtobits(-0.1463422),$shortrealtobits(-0.060737316),$shortrealtobits(-0.35839006),
    $shortrealtobits(-0.23079027),$shortrealtobits(0.28280434),$shortrealtobits(-0.47914347),$shortrealtobits(0.22066016),
    $shortrealtobits(-0.13891014),$shortrealtobits(-0.46581483),$shortrealtobits(-0.31236172),$shortrealtobits(0.5795618),
    $shortrealtobits(0.12867585),$shortrealtobits(-0.33881167),$shortrealtobits(0.35092965),$shortrealtobits(-0.46622577),
    $shortrealtobits(-0.25764737),$shortrealtobits(0.30567965),$shortrealtobits(0.30329472),$shortrealtobits(-0.4926346)
  },
  '{ 
    $shortrealtobits(0.014531706),$shortrealtobits(0.43891257),$shortrealtobits(-0.0068248585),$shortrealtobits(0.061848048),
    $shortrealtobits(0.34919152),$shortrealtobits(0.38228732),$shortrealtobits(-0.2745033),$shortrealtobits(0.0013365367),
    $shortrealtobits(0.1677584),$shortrealtobits(0.4001345),$shortrealtobits(0.37049094),$shortrealtobits(0.11412082),
    $shortrealtobits(0.27424285),$shortrealtobits(-0.2531464),$shortrealtobits(0.2649959),$shortrealtobits(0.4379082),
    $shortrealtobits(0.16071273),$shortrealtobits(0.10520196),$shortrealtobits(-0.07190809),$shortrealtobits(-0.18150018),
    $shortrealtobits(0.4598873),$shortrealtobits(-0.023676293),$shortrealtobits(-0.054034986),$shortrealtobits(0.17654963),
    $shortrealtobits(0.15859531),$shortrealtobits(0.4639537),$shortrealtobits(-0.26229417),$shortrealtobits(-0.34869555),
    $shortrealtobits(-0.030834908),$shortrealtobits(-0.11662379),$shortrealtobits(0.13794635),$shortrealtobits(-0.15588304),
    $shortrealtobits(0.4316786),$shortrealtobits(-0.3510806),$shortrealtobits(0.11240149),$shortrealtobits(0.18208055),
    $shortrealtobits(0.2233249),$shortrealtobits(0.024962487),$shortrealtobits(-0.21023957),$shortrealtobits(-0.083141916)
  },
  '{ 
    $shortrealtobits(0.6922004),$shortrealtobits(0.025198488),$shortrealtobits(0.34569314),$shortrealtobits(0.44642535),
    $shortrealtobits(-0.28739226),$shortrealtobits(-0.121381484),$shortrealtobits(-0.30677196),$shortrealtobits(-0.3006623),
    $shortrealtobits(0.4219753),$shortrealtobits(0.39431414),$shortrealtobits(0.018517552),$shortrealtobits(-0.44955218),
    $shortrealtobits(-0.075195245),$shortrealtobits(0.052924145),$shortrealtobits(-0.19784),$shortrealtobits(0.24436177),
    $shortrealtobits(-0.027502075),$shortrealtobits(0.07088162),$shortrealtobits(0.15332958),$shortrealtobits(0.0990803),
    $shortrealtobits(-0.10154435),$shortrealtobits(0.30637527),$shortrealtobits(-0.003215529),$shortrealtobits(0.103054546),
    $shortrealtobits(0.29098058),$shortrealtobits(-0.23515573),$shortrealtobits(-0.19617589),$shortrealtobits(-0.68993497),
    $shortrealtobits(-0.22641668),$shortrealtobits(0.13568017),$shortrealtobits(-0.48904023),$shortrealtobits(-0.6765585),
    $shortrealtobits(0.25893185),$shortrealtobits(0.14702733),$shortrealtobits(0.09226928),$shortrealtobits(-0.09695095),
    $shortrealtobits(0.23526111),$shortrealtobits(-0.24489239),$shortrealtobits(-0.24931398),$shortrealtobits(-0.046659324)
  },
  '{ 
    $shortrealtobits(0.5521156),$shortrealtobits(-0.25635353),$shortrealtobits(-0.0626214),$shortrealtobits(-0.46526656),
    $shortrealtobits(0.30999586),$shortrealtobits(-0.17965595),$shortrealtobits(0.12422267),$shortrealtobits(-0.38124517),
    $shortrealtobits(0.42349097),$shortrealtobits(0.830878),$shortrealtobits(-0.46300325),$shortrealtobits(-0.12994741),
    $shortrealtobits(-0.1430227),$shortrealtobits(0.13847466),$shortrealtobits(0.10234797),$shortrealtobits(-0.15857835),
    $shortrealtobits(0.53010553),$shortrealtobits(-0.021374037),$shortrealtobits(-0.08302116),$shortrealtobits(-0.104123674),
    $shortrealtobits(0.21032052),$shortrealtobits(0.060323983),$shortrealtobits(-0.2291589),$shortrealtobits(-0.2153842),
    $shortrealtobits(-0.017616812),$shortrealtobits(-0.2876413),$shortrealtobits(0.3482484),$shortrealtobits(0.33218443),
    $shortrealtobits(-0.2324995),$shortrealtobits(0.106761046),$shortrealtobits(0.3595252),$shortrealtobits(-0.3542829),
    $shortrealtobits(0.056635525),$shortrealtobits(-0.4759693),$shortrealtobits(0.6435635),$shortrealtobits(-0.0790747),
    $shortrealtobits(0.17766528),$shortrealtobits(-0.004368377),$shortrealtobits(-0.21677119),$shortrealtobits(0.34683025)
  },
  '{ 
    $shortrealtobits(0.15518805),$shortrealtobits(-0.33325264),$shortrealtobits(-0.42067838),$shortrealtobits(0.37264392),
    $shortrealtobits(0.033477966),$shortrealtobits(-0.27378273),$shortrealtobits(0.44956443),$shortrealtobits(0.033890173),
    $shortrealtobits(0.3619253),$shortrealtobits(-0.47859457),$shortrealtobits(-0.06996032),$shortrealtobits(0.46401227),
    $shortrealtobits(0.3559901),$shortrealtobits(0.36069328),$shortrealtobits(-0.33233163),$shortrealtobits(-0.32411137),
    $shortrealtobits(-0.75999534),$shortrealtobits(0.28742886),$shortrealtobits(-0.022140551),$shortrealtobits(0.09123756),
    $shortrealtobits(-0.05341973),$shortrealtobits(-0.42007306),$shortrealtobits(-0.47674444),$shortrealtobits(-0.40057653),
    $shortrealtobits(-0.17885849),$shortrealtobits(0.08838895),$shortrealtobits(-0.2908125),$shortrealtobits(-0.1046324),
    $shortrealtobits(0.48373342),$shortrealtobits(-0.021994276),$shortrealtobits(-0.0071373773),$shortrealtobits(0.33331746),
    $shortrealtobits(0.35478652),$shortrealtobits(-0.022076698),$shortrealtobits(-0.045248084),$shortrealtobits(0.095024206),
    $shortrealtobits(0.42158073),$shortrealtobits(0.38794068),$shortrealtobits(0.08629065),$shortrealtobits(-0.08484484)
  },
  '{ 
    $shortrealtobits(0.06528808),$shortrealtobits(-0.16758868),$shortrealtobits(-0.15223527),$shortrealtobits(0.044104766),
    $shortrealtobits(-0.003917477),$shortrealtobits(-0.13900065),$shortrealtobits(-0.013663963),$shortrealtobits(0.35793754),
    $shortrealtobits(-0.17168887),$shortrealtobits(-0.23014842),$shortrealtobits(0.27622876),$shortrealtobits(0.01009628),
    $shortrealtobits(-0.009280202),$shortrealtobits(-0.20003842),$shortrealtobits(0.07504048),$shortrealtobits(0.3383062),
    $shortrealtobits(-0.44532135),$shortrealtobits(0.26206088),$shortrealtobits(-0.06080208),$shortrealtobits(-0.54262257),
    $shortrealtobits(0.3053301),$shortrealtobits(0.053276274),$shortrealtobits(0.08583672),$shortrealtobits(-0.20106879),
    $shortrealtobits(0.33830726),$shortrealtobits(0.47461057),$shortrealtobits(-0.6327542),$shortrealtobits(-0.11135385),
    $shortrealtobits(-0.05642195),$shortrealtobits(0.07744964),$shortrealtobits(-0.2942699),$shortrealtobits(-0.4011981),
    $shortrealtobits(0.10448533),$shortrealtobits(-0.056507017),$shortrealtobits(0.030613633),$shortrealtobits(0.10167322),
    $shortrealtobits(-0.23172125),$shortrealtobits(-0.25394726),$shortrealtobits(-0.31323594),$shortrealtobits(-0.22560014)
  },
  '{ 
    $shortrealtobits(-0.0029893708),$shortrealtobits(0.39705244),$shortrealtobits(-0.23851232),$shortrealtobits(0.23255062),
    $shortrealtobits(0.6058438),$shortrealtobits(0.23459126),$shortrealtobits(0.24567273),$shortrealtobits(0.35098237),
    $shortrealtobits(-0.12699981),$shortrealtobits(0.1577117),$shortrealtobits(0.0080418065),$shortrealtobits(-0.3323296),
    $shortrealtobits(-0.0428255),$shortrealtobits(0.492639),$shortrealtobits(0.4003864),$shortrealtobits(0.45155975),
    $shortrealtobits(-0.09912736),$shortrealtobits(-0.014794579),$shortrealtobits(-0.07669835),$shortrealtobits(-0.025018847),
    $shortrealtobits(0.12148393),$shortrealtobits(0.31271225),$shortrealtobits(-0.0052804984),$shortrealtobits(0.0715828),
    $shortrealtobits(-0.46121395),$shortrealtobits(0.24281545),$shortrealtobits(0.39294058),$shortrealtobits(-0.052655693),
    $shortrealtobits(0.39723164),$shortrealtobits(-0.10481112),$shortrealtobits(0.35389072),$shortrealtobits(0.3318103),
    $shortrealtobits(-0.27156353),$shortrealtobits(0.119682655),$shortrealtobits(-0.14679512),$shortrealtobits(0.11947784),
    $shortrealtobits(-0.079209894),$shortrealtobits(-0.049740095),$shortrealtobits(0.32665566),$shortrealtobits(0.24363378)
  },
  '{ 
    $shortrealtobits(-0.018619802),$shortrealtobits(0.22412032),$shortrealtobits(0.1655088),$shortrealtobits(-0.48055702),
    $shortrealtobits(0.21744832),$shortrealtobits(-0.39709052),$shortrealtobits(-0.36781123),$shortrealtobits(0.62694293),
    $shortrealtobits(0.22675553),$shortrealtobits(0.042914975),$shortrealtobits(0.38321057),$shortrealtobits(-0.1539923),
    $shortrealtobits(0.04345159),$shortrealtobits(-0.09145994),$shortrealtobits(0.02191905),$shortrealtobits(0.35804313),
    $shortrealtobits(0.31548604),$shortrealtobits(0.07160174),$shortrealtobits(0.32748073),$shortrealtobits(-0.5289925),
    $shortrealtobits(-0.38047937),$shortrealtobits(0.4057355),$shortrealtobits(0.21219008),$shortrealtobits(0.06707627),
    $shortrealtobits(0.02512561),$shortrealtobits(0.2895732),$shortrealtobits(-0.5679257),$shortrealtobits(0.10964277),
    $shortrealtobits(-0.35698712),$shortrealtobits(0.3681122),$shortrealtobits(0.11214821),$shortrealtobits(-0.41201043),
    $shortrealtobits(0.22340606),$shortrealtobits(-0.46108487),$shortrealtobits(-0.14752412),$shortrealtobits(0.31994727),
    $shortrealtobits(0.14709158),$shortrealtobits(0.11651058),$shortrealtobits(0.38611442),$shortrealtobits(-0.38168585)
  },
  '{ 
    $shortrealtobits(-0.069771945),$shortrealtobits(-0.3808906),$shortrealtobits(-0.04816783),$shortrealtobits(-0.24956805),
    $shortrealtobits(0.27330574),$shortrealtobits(-0.4723528),$shortrealtobits(0.49032637),$shortrealtobits(-0.06920525),
    $shortrealtobits(-0.45816278),$shortrealtobits(0.39580032),$shortrealtobits(-0.113338284),$shortrealtobits(0.530343),
    $shortrealtobits(-0.099556446),$shortrealtobits(-0.10972891),$shortrealtobits(0.4693019),$shortrealtobits(0.20458671),
    $shortrealtobits(-0.36835986),$shortrealtobits(0.7216057),$shortrealtobits(-0.27180487),$shortrealtobits(-0.33355436),
    $shortrealtobits(0.25989535),$shortrealtobits(0.30792162),$shortrealtobits(0.028868355),$shortrealtobits(0.3329948),
    $shortrealtobits(-0.18883674),$shortrealtobits(-0.12043692),$shortrealtobits(-0.5954286),$shortrealtobits(0.5800862),
    $shortrealtobits(-0.59340274),$shortrealtobits(0.37300277),$shortrealtobits(0.24245362),$shortrealtobits(-0.3484739),
    $shortrealtobits(0.33017886),$shortrealtobits(0.22705899),$shortrealtobits(0.05426448),$shortrealtobits(-0.059487224),
    $shortrealtobits(0.4302596),$shortrealtobits(-0.29526073),$shortrealtobits(0.23638274),$shortrealtobits(-0.51894724)
  },
  '{ 
    $shortrealtobits(0.03131434),$shortrealtobits(-0.14521608),$shortrealtobits(0.32874548),$shortrealtobits(0.3432401),
    $shortrealtobits(-0.35737565),$shortrealtobits(-0.7160062),$shortrealtobits(0.11964594),$shortrealtobits(-0.28769645),
    $shortrealtobits(-0.5645043),$shortrealtobits(0.20861247),$shortrealtobits(0.754159),$shortrealtobits(-0.36944288),
    $shortrealtobits(0.11333746),$shortrealtobits(0.5120868),$shortrealtobits(-0.59111696),$shortrealtobits(-0.08572931),
    $shortrealtobits(-0.23645489),$shortrealtobits(-0.07999221),$shortrealtobits(0.2198535),$shortrealtobits(-0.48670873),
    $shortrealtobits(0.016465703),$shortrealtobits(0.24303837),$shortrealtobits(0.06484045),$shortrealtobits(0.4480264),
    $shortrealtobits(0.22207156),$shortrealtobits(0.2015675),$shortrealtobits(0.31782588),$shortrealtobits(0.12091812),
    $shortrealtobits(0.24195823),$shortrealtobits(-0.46246958),$shortrealtobits(0.40213993),$shortrealtobits(-0.024512252),
    $shortrealtobits(0.43799627),$shortrealtobits(-0.22373325),$shortrealtobits(-0.046105094),$shortrealtobits(0.28352642),
    $shortrealtobits(0.303697),$shortrealtobits(0.08545675),$shortrealtobits(-0.043038722),$shortrealtobits(0.28182593)
  },
  '{ 
    $shortrealtobits(-0.36412144),$shortrealtobits(0.19816709),$shortrealtobits(0.2609341),$shortrealtobits(0.21026455),
    $shortrealtobits(0.1765886),$shortrealtobits(0.0022401356),$shortrealtobits(0.8023658),$shortrealtobits(0.27152893),
    $shortrealtobits(0.22701406),$shortrealtobits(0.0130867055),$shortrealtobits(-0.025584199),$shortrealtobits(0.4490657),
    $shortrealtobits(0.1638749),$shortrealtobits(0.44304702),$shortrealtobits(-0.42099333),$shortrealtobits(-0.13485695),
    $shortrealtobits(-0.118206926),$shortrealtobits(-0.17231324),$shortrealtobits(-0.14566827),$shortrealtobits(0.4171778),
    $shortrealtobits(-0.4579135),$shortrealtobits(0.2207391),$shortrealtobits(0.33172166),$shortrealtobits(-0.49229896),
    $shortrealtobits(-0.13967274),$shortrealtobits(-0.014978187),$shortrealtobits(0.6039107),$shortrealtobits(-0.71133286),
    $shortrealtobits(0.6939044),$shortrealtobits(-0.13692105),$shortrealtobits(-0.30777857),$shortrealtobits(-0.7340108),
    $shortrealtobits(-0.34641114),$shortrealtobits(0.12791722),$shortrealtobits(0.26996338),$shortrealtobits(0.48154762),
    $shortrealtobits(0.24211827),$shortrealtobits(0.17744143),$shortrealtobits(0.037961584),$shortrealtobits(0.63231254)
  },
  '{ 
    $shortrealtobits(0.6177302),$shortrealtobits(-0.19420838),$shortrealtobits(-0.19028705),$shortrealtobits(-0.044989105),
    $shortrealtobits(-0.22304444),$shortrealtobits(0.5406044),$shortrealtobits(0.32207957),$shortrealtobits(-0.40143698),
    $shortrealtobits(-0.1960274),$shortrealtobits(-0.3549164),$shortrealtobits(0.19858335),$shortrealtobits(0.038842164),
    $shortrealtobits(-0.0046261935),$shortrealtobits(-0.29020742),$shortrealtobits(-0.37473923),$shortrealtobits(-0.3826141),
    $shortrealtobits(-0.5486989),$shortrealtobits(-0.54534173),$shortrealtobits(-0.110318206),$shortrealtobits(0.46570632),
    $shortrealtobits(-0.14627677),$shortrealtobits(0.26396906),$shortrealtobits(0.4564492),$shortrealtobits(-0.31299415),
    $shortrealtobits(0.012002592),$shortrealtobits(-0.45239112),$shortrealtobits(-0.6888782),$shortrealtobits(-0.33480737),
    $shortrealtobits(-0.17955261),$shortrealtobits(-0.07972104),$shortrealtobits(-0.16931196),$shortrealtobits(-0.0068548955),
    $shortrealtobits(-0.38668936),$shortrealtobits(-0.37721542),$shortrealtobits(0.17908777),$shortrealtobits(0.16555665),
    $shortrealtobits(0.28345838),$shortrealtobits(-0.41105768),$shortrealtobits(-0.16471335),$shortrealtobits(-0.2895481)
  },
  '{ 
    $shortrealtobits(0.21894395),$shortrealtobits(-0.36440802),$shortrealtobits(-0.12463689),$shortrealtobits(-0.33165297),
    $shortrealtobits(-0.019305699),$shortrealtobits(-0.31331468),$shortrealtobits(-0.3159665),$shortrealtobits(-0.4146383),
    $shortrealtobits(-0.26229966),$shortrealtobits(0.42133147),$shortrealtobits(0.2509268),$shortrealtobits(-0.30946964),
    $shortrealtobits(-0.25395665),$shortrealtobits(0.42841753),$shortrealtobits(0.16009296),$shortrealtobits(0.15080711),
    $shortrealtobits(0.2914993),$shortrealtobits(0.39713928),$shortrealtobits(-0.26259127),$shortrealtobits(0.13405411),
    $shortrealtobits(0.12066404),$shortrealtobits(0.11376942),$shortrealtobits(0.43128082),$shortrealtobits(0.4548441),
    $shortrealtobits(0.12258066),$shortrealtobits(0.05541075),$shortrealtobits(0.020574534),$shortrealtobits(-0.34894603),
    $shortrealtobits(-0.42359188),$shortrealtobits(0.17906147),$shortrealtobits(0.5425973),$shortrealtobits(-0.08653047),
    $shortrealtobits(-0.4764079),$shortrealtobits(0.37033823),$shortrealtobits(0.19284703),$shortrealtobits(-0.17607935),
    $shortrealtobits(0.47518492),$shortrealtobits(-0.42511234),$shortrealtobits(-0.45368955),$shortrealtobits(0.022263845)
  },
  '{ 
    $shortrealtobits(-0.63389444),$shortrealtobits(-0.5333558),$shortrealtobits(0.26418316),$shortrealtobits(-0.3098004),
    $shortrealtobits(-0.2863051),$shortrealtobits(0.22391209),$shortrealtobits(-0.1549494),$shortrealtobits(0.14211282),
    $shortrealtobits(-0.6066439),$shortrealtobits(0.028001653),$shortrealtobits(-0.5113389),$shortrealtobits(0.16962983),
    $shortrealtobits(0.04898956),$shortrealtobits(0.09056523),$shortrealtobits(-0.35826176),$shortrealtobits(0.06491407),
    $shortrealtobits(0.23268653),$shortrealtobits(-0.085400894),$shortrealtobits(-0.42297444),$shortrealtobits(0.38841945),
    $shortrealtobits(0.24319297),$shortrealtobits(-0.30387765),$shortrealtobits(-0.5993262),$shortrealtobits(0.3103772),
    $shortrealtobits(-0.30987623),$shortrealtobits(0.510765),$shortrealtobits(-0.3539893),$shortrealtobits(-0.081063144),
    $shortrealtobits(0.6599169),$shortrealtobits(-0.28341603),$shortrealtobits(-0.2225057),$shortrealtobits(-0.17991005),
    $shortrealtobits(0.2516483),$shortrealtobits(-0.014039973),$shortrealtobits(-0.2844877),$shortrealtobits(0.41843095),
    $shortrealtobits(-0.15106738),$shortrealtobits(-0.14356162),$shortrealtobits(-0.4588769),$shortrealtobits(0.07059036)
  },
  '{ 
    $shortrealtobits(-0.25558555),$shortrealtobits(0.12119865),$shortrealtobits(-0.42199045),$shortrealtobits(-0.1831091),
    $shortrealtobits(-0.13345674),$shortrealtobits(0.24072537),$shortrealtobits(0.10084306),$shortrealtobits(0.36008817),
    $shortrealtobits(0.31555626),$shortrealtobits(-0.26922363),$shortrealtobits(0.6243971),$shortrealtobits(-0.13202848),
    $shortrealtobits(-0.38921434),$shortrealtobits(-0.2935741),$shortrealtobits(-0.36321324),$shortrealtobits(0.56765693),
    $shortrealtobits(0.3834301),$shortrealtobits(0.10289531),$shortrealtobits(-0.39086556),$shortrealtobits(-0.20743692),
    $shortrealtobits(-0.539165),$shortrealtobits(-0.03639045),$shortrealtobits(-0.46916336),$shortrealtobits(0.18767907),
    $shortrealtobits(-0.24497956),$shortrealtobits(0.4523702),$shortrealtobits(-0.13159166),$shortrealtobits(0.059371646),
    $shortrealtobits(-0.27333173),$shortrealtobits(-0.4755338),$shortrealtobits(-0.075812235),$shortrealtobits(0.31860033),
    $shortrealtobits(0.47097683),$shortrealtobits(-0.46233925),$shortrealtobits(-0.010709581),$shortrealtobits(0.207593),
    $shortrealtobits(-0.31345856),$shortrealtobits(-0.04392105),$shortrealtobits(0.63565147),$shortrealtobits(0.07157847)
  },
  '{ 
    $shortrealtobits(-0.011406712),$shortrealtobits(-0.13954443),$shortrealtobits(-0.50957656),$shortrealtobits(0.27780604),
    $shortrealtobits(0.71297556),$shortrealtobits(0.0034561579),$shortrealtobits(-0.032380942),$shortrealtobits(-0.00090557226),
    $shortrealtobits(0.14833885),$shortrealtobits(0.18090612),$shortrealtobits(-0.8343409),$shortrealtobits(0.18592194),
    $shortrealtobits(-0.31902683),$shortrealtobits(-0.30555344),$shortrealtobits(0.35316542),$shortrealtobits(-0.37376294),
    $shortrealtobits(0.18590714),$shortrealtobits(-0.032531444),$shortrealtobits(-0.058240443),$shortrealtobits(-0.07621346),
    $shortrealtobits(-0.15069725),$shortrealtobits(-0.23045076),$shortrealtobits(0.37356174),$shortrealtobits(-0.08178507),
    $shortrealtobits(0.24004327),$shortrealtobits(0.2897285),$shortrealtobits(-0.1989463),$shortrealtobits(0.4069787),
    $shortrealtobits(0.021354945),$shortrealtobits(-0.5497931),$shortrealtobits(-0.05930171),$shortrealtobits(0.6015351),
    $shortrealtobits(-0.490338),$shortrealtobits(-0.3605671),$shortrealtobits(-0.1761273),$shortrealtobits(-0.03439894),
    $shortrealtobits(0.27383688),$shortrealtobits(-0.13612017),$shortrealtobits(0.03993376),$shortrealtobits(-0.26352093)
  },
  '{ 
    $shortrealtobits(-0.19305354),$shortrealtobits(0.6269849),$shortrealtobits(0.12373783),$shortrealtobits(0.20858651),
    $shortrealtobits(-0.12439302),$shortrealtobits(0.017745959),$shortrealtobits(-0.17461462),$shortrealtobits(-0.124870114),
    $shortrealtobits(0.14902271),$shortrealtobits(-0.13172098),$shortrealtobits(-0.04390849),$shortrealtobits(-0.38467738),
    $shortrealtobits(0.2054493),$shortrealtobits(0.10448262),$shortrealtobits(-0.38497913),$shortrealtobits(0.25677523),
    $shortrealtobits(0.3792274),$shortrealtobits(0.17755641),$shortrealtobits(0.13486134),$shortrealtobits(-0.20767732),
    $shortrealtobits(0.16107279),$shortrealtobits(-0.20824277),$shortrealtobits(-0.3147227),$shortrealtobits(-0.4364213),
    $shortrealtobits(0.24678423),$shortrealtobits(0.24935108),$shortrealtobits(-0.03329508),$shortrealtobits(0.41967285),
    $shortrealtobits(-0.5845927),$shortrealtobits(-0.38139483),$shortrealtobits(0.31991923),$shortrealtobits(0.6779165),
    $shortrealtobits(-0.30527782),$shortrealtobits(0.19282915),$shortrealtobits(0.18281688),$shortrealtobits(-0.2909022),
    $shortrealtobits(0.54246664),$shortrealtobits(0.22550547),$shortrealtobits(0.31782973),$shortrealtobits(0.023550272)
  },
  '{ 
    $shortrealtobits(-0.21879952),$shortrealtobits(0.094545856),$shortrealtobits(0.053476155),$shortrealtobits(0.029741375),
    $shortrealtobits(-0.2612455),$shortrealtobits(-0.10480306),$shortrealtobits(-0.23806182),$shortrealtobits(-0.3068835),
    $shortrealtobits(-0.13424173),$shortrealtobits(0.0055004456),$shortrealtobits(-0.066339776),$shortrealtobits(0.26279965),
    $shortrealtobits(0.31052586),$shortrealtobits(0.037678085),$shortrealtobits(0.23232703),$shortrealtobits(-0.30992252),
    $shortrealtobits(0.26921156),$shortrealtobits(0.1871889),$shortrealtobits(0.44545886),$shortrealtobits(0.014562807),
    $shortrealtobits(-0.36426106),$shortrealtobits(0.16105358),$shortrealtobits(0.031086454),$shortrealtobits(0.9891883),
    $shortrealtobits(-0.32665482),$shortrealtobits(0.39432418),$shortrealtobits(-0.6467474),$shortrealtobits(-0.6690666),
    $shortrealtobits(0.46747395),$shortrealtobits(-0.4279193),$shortrealtobits(-0.35424906),$shortrealtobits(0.25718036),
    $shortrealtobits(0.37312007),$shortrealtobits(0.26989844),$shortrealtobits(-0.6892061),$shortrealtobits(0.5282656),
    $shortrealtobits(-0.066132665),$shortrealtobits(-0.013296257),$shortrealtobits(0.06924483),$shortrealtobits(-0.66906375)
  },
  '{ 
    $shortrealtobits(0.17978865),$shortrealtobits(0.18067048),$shortrealtobits(0.117577486),$shortrealtobits(0.090568535),
    $shortrealtobits(-0.5280929),$shortrealtobits(-0.2063946),$shortrealtobits(-0.75201553),$shortrealtobits(-0.46872842),
    $shortrealtobits(0.15234509),$shortrealtobits(0.10423144),$shortrealtobits(0.25711775),$shortrealtobits(-0.34741998),
    $shortrealtobits(-0.1871383),$shortrealtobits(0.097559825),$shortrealtobits(0.06914299),$shortrealtobits(0.050983503),
    $shortrealtobits(-0.17298093),$shortrealtobits(-0.023039343),$shortrealtobits(-0.38230792),$shortrealtobits(0.6101223),
    $shortrealtobits(0.46083924),$shortrealtobits(0.19794223),$shortrealtobits(0.18504325),$shortrealtobits(0.022318263),
    $shortrealtobits(0.41026422),$shortrealtobits(0.15504774),$shortrealtobits(-0.04036512),$shortrealtobits(-0.30813816),
    $shortrealtobits(-0.18692872),$shortrealtobits(0.095282964),$shortrealtobits(0.6287247),$shortrealtobits(0.06986608),
    $shortrealtobits(0.22831164),$shortrealtobits(-0.4457293),$shortrealtobits(0.11829689),$shortrealtobits(-0.38473263),
    $shortrealtobits(-0.3281319),$shortrealtobits(0.22250775),$shortrealtobits(-0.31146067),$shortrealtobits(-0.5959563)
  },
  '{ 
    $shortrealtobits(0.8745724),$shortrealtobits(0.101702094),$shortrealtobits(0.7325185),$shortrealtobits(-0.11540211),
    $shortrealtobits(-0.06804807),$shortrealtobits(-0.06830655),$shortrealtobits(-0.32350025),$shortrealtobits(-0.13723461),
    $shortrealtobits(0.17455623),$shortrealtobits(-0.24909149),$shortrealtobits(0.2273687),$shortrealtobits(0.28331757),
    $shortrealtobits(-0.24169838),$shortrealtobits(-0.41910747),$shortrealtobits(0.2096112),$shortrealtobits(0.12046535),
    $shortrealtobits(-0.17045696),$shortrealtobits(-0.335277),$shortrealtobits(-0.25111955),$shortrealtobits(-0.06445309),
    $shortrealtobits(0.1579041),$shortrealtobits(0.3993323),$shortrealtobits(0.21889365),$shortrealtobits(-0.38077983),
    $shortrealtobits(-0.00899804),$shortrealtobits(0.28863487),$shortrealtobits(-0.1292636),$shortrealtobits(-0.09559274),
    $shortrealtobits(0.041669793),$shortrealtobits(0.0030956396),$shortrealtobits(0.112000085),$shortrealtobits(0.23149861),
    $shortrealtobits(0.020190531),$shortrealtobits(-0.0019297258),$shortrealtobits(0.05941593),$shortrealtobits(0.21795052),
    $shortrealtobits(-0.2367467),$shortrealtobits(-0.22677822),$shortrealtobits(0.27120385),$shortrealtobits(0.29189056)
  },
  '{ 
    $shortrealtobits(0.20640719),$shortrealtobits(-0.11139871),$shortrealtobits(0.71547747),$shortrealtobits(0.49441016),
    $shortrealtobits(0.12325753),$shortrealtobits(0.09848645),$shortrealtobits(0.024023192),$shortrealtobits(-0.36001077),
    $shortrealtobits(-0.40893677),$shortrealtobits(-0.34161216),$shortrealtobits(-0.16103524),$shortrealtobits(-0.08648441),
    $shortrealtobits(0.2716748),$shortrealtobits(0.11139701),$shortrealtobits(-0.4682231),$shortrealtobits(-0.25740337),
    $shortrealtobits(-0.35516074),$shortrealtobits(0.35220525),$shortrealtobits(0.11605947),$shortrealtobits(0.36086127),
    $shortrealtobits(0.005561749),$shortrealtobits(-0.020675216),$shortrealtobits(0.49014977),$shortrealtobits(-0.28385046),
    $shortrealtobits(0.4405696),$shortrealtobits(-0.4690474),$shortrealtobits(0.33035898),$shortrealtobits(0.08510705),
    $shortrealtobits(0.24533255),$shortrealtobits(-0.054696836),$shortrealtobits(0.14501494),$shortrealtobits(-0.10894127),
    $shortrealtobits(0.15240136),$shortrealtobits(-0.08931054),$shortrealtobits(0.16484748),$shortrealtobits(0.2546626),
    $shortrealtobits(0.09398579),$shortrealtobits(-0.2736664),$shortrealtobits(-0.24326305),$shortrealtobits(0.47175112)
  },
  '{ 
    $shortrealtobits(0.010980269),$shortrealtobits(-0.21871553),$shortrealtobits(0.046689723),$shortrealtobits(0.4942887),
    $shortrealtobits(0.26265538),$shortrealtobits(-0.10949712),$shortrealtobits(0.21501821),$shortrealtobits(-0.28028774),
    $shortrealtobits(-0.40322742),$shortrealtobits(-0.38415122),$shortrealtobits(-0.03294176),$shortrealtobits(-0.17735498),
    $shortrealtobits(0.16018365),$shortrealtobits(-0.02044588),$shortrealtobits(-0.2709275),$shortrealtobits(-0.35246995),
    $shortrealtobits(0.28638327),$shortrealtobits(0.46494788),$shortrealtobits(-0.112465516),$shortrealtobits(-0.1498194),
    $shortrealtobits(0.19193451),$shortrealtobits(0.5592275),$shortrealtobits(0.1702718),$shortrealtobits(0.03415536),
    $shortrealtobits(0.12152552),$shortrealtobits(0.28639108),$shortrealtobits(-0.033794977),$shortrealtobits(-0.19356768),
    $shortrealtobits(-0.3867313),$shortrealtobits(0.095718),$shortrealtobits(0.39038715),$shortrealtobits(-0.48290294),
    $shortrealtobits(0.090904236),$shortrealtobits(0.55224776),$shortrealtobits(0.62177074),$shortrealtobits(-0.26892778),
    $shortrealtobits(-0.25698894),$shortrealtobits(0.515741),$shortrealtobits(-0.12956485),$shortrealtobits(0.16559365)
  },
  '{ 
    $shortrealtobits(-0.0464036),$shortrealtobits(0.41032863),$shortrealtobits(-0.20040193),$shortrealtobits(-0.16781835),
    $shortrealtobits(-0.46486852),$shortrealtobits(-0.32225397),$shortrealtobits(0.40928632),$shortrealtobits(-0.20821133),
    $shortrealtobits(-0.1267124),$shortrealtobits(-0.24706984),$shortrealtobits(-0.27782923),$shortrealtobits(0.1668109),
    $shortrealtobits(0.24288926),$shortrealtobits(-0.42441964),$shortrealtobits(-0.11941708),$shortrealtobits(-0.19737367),
    $shortrealtobits(0.14717568),$shortrealtobits(0.042132713),$shortrealtobits(0.55149716),$shortrealtobits(-0.018714914),
    $shortrealtobits(-0.41087258),$shortrealtobits(0.29089448),$shortrealtobits(0.305439),$shortrealtobits(-0.38556033),
    $shortrealtobits(0.08911588),$shortrealtobits(-0.28859648),$shortrealtobits(0.39094526),$shortrealtobits(-0.29657224),
    $shortrealtobits(-0.026131734),$shortrealtobits(0.35330942),$shortrealtobits(0.2938475),$shortrealtobits(-0.31873786),
    $shortrealtobits(-0.1774912),$shortrealtobits(0.40001947),$shortrealtobits(0.45131832),$shortrealtobits(-0.050962925),
    $shortrealtobits(0.23914339),$shortrealtobits(0.2549366),$shortrealtobits(0.4633777),$shortrealtobits(-0.026163863)
  },
  '{ 
    $shortrealtobits(-0.47465762),$shortrealtobits(0.30179504),$shortrealtobits(-0.23516186),$shortrealtobits(0.16052426),
    $shortrealtobits(0.14510687),$shortrealtobits(-0.14917059),$shortrealtobits(0.003989333),$shortrealtobits(-0.21895002),
    $shortrealtobits(-0.15822783),$shortrealtobits(0.35957807),$shortrealtobits(-0.039243013),$shortrealtobits(-0.27145827),
    $shortrealtobits(-0.16938676),$shortrealtobits(-0.009496244),$shortrealtobits(0.18642034),$shortrealtobits(0.024455853),
    $shortrealtobits(-0.10308975),$shortrealtobits(-0.103707746),$shortrealtobits(-0.1465259),$shortrealtobits(-0.12663674),
    $shortrealtobits(0.33081976),$shortrealtobits(0.22281955),$shortrealtobits(-0.33043906),$shortrealtobits(0.3554844),
    $shortrealtobits(0.35226774),$shortrealtobits(-0.13904463),$shortrealtobits(-0.39581573),$shortrealtobits(-0.26789203),
    $shortrealtobits(-0.044651918),$shortrealtobits(0.107426256),$shortrealtobits(-0.12772366),$shortrealtobits(-0.0925649),
    $shortrealtobits(-0.50357264),$shortrealtobits(0.10630806),$shortrealtobits(-0.22240475),$shortrealtobits(0.14765814),
    $shortrealtobits(0.07122923),$shortrealtobits(0.48014116),$shortrealtobits(-0.30219105),$shortrealtobits(0.09276434)
  },
  '{ 
    $shortrealtobits(0.42151865),$shortrealtobits(-0.8170706),$shortrealtobits(-0.015640343),$shortrealtobits(-0.45911345),
    $shortrealtobits(0.06471275),$shortrealtobits(0.0048445635),$shortrealtobits(-0.1783796),$shortrealtobits(-0.20214437),
    $shortrealtobits(0.32825285),$shortrealtobits(0.07946046),$shortrealtobits(-0.4401781),$shortrealtobits(0.41854084),
    $shortrealtobits(-0.11073019),$shortrealtobits(-0.050461374),$shortrealtobits(-0.4096857),$shortrealtobits(0.18941516),
    $shortrealtobits(-0.31264034),$shortrealtobits(-0.16616471),$shortrealtobits(-0.048044186),$shortrealtobits(-0.14945713),
    $shortrealtobits(-0.22501305),$shortrealtobits(-0.44135818),$shortrealtobits(0.41770032),$shortrealtobits(0.07130177),
    $shortrealtobits(0.24663061),$shortrealtobits(-0.044959333),$shortrealtobits(0.28662792),$shortrealtobits(0.17808194),
    $shortrealtobits(0.027140463),$shortrealtobits(0.23782405),$shortrealtobits(-0.030443914),$shortrealtobits(0.21831575),
    $shortrealtobits(-0.40153256),$shortrealtobits(-0.337079),$shortrealtobits(-0.2639012),$shortrealtobits(0.39710304),
    $shortrealtobits(0.19788393),$shortrealtobits(-0.3066279),$shortrealtobits(0.23884757),$shortrealtobits(-0.042075284)
  },
  '{ 
    $shortrealtobits(0.20448467),$shortrealtobits(0.21316889),$shortrealtobits(-0.32037148),$shortrealtobits(0.096687935),
    $shortrealtobits(0.28682154),$shortrealtobits(-0.43043143),$shortrealtobits(0.6480322),$shortrealtobits(0.46653625),
    $shortrealtobits(-0.32588506),$shortrealtobits(-0.019104516),$shortrealtobits(0.4320713),$shortrealtobits(0.5240076),
    $shortrealtobits(-0.55449957),$shortrealtobits(-0.07434075),$shortrealtobits(0.4337765),$shortrealtobits(0.5204722),
    $shortrealtobits(0.2434616),$shortrealtobits(0.18203028),$shortrealtobits(-0.43354443),$shortrealtobits(-0.5382657),
    $shortrealtobits(0.17689858),$shortrealtobits(0.010938741),$shortrealtobits(0.31443256),$shortrealtobits(-0.38983262),
    $shortrealtobits(0.16561146),$shortrealtobits(0.5323758),$shortrealtobits(0.46329483),$shortrealtobits(-0.2382617),
    $shortrealtobits(0.4979657),$shortrealtobits(0.24994655),$shortrealtobits(-0.031569973),$shortrealtobits(-0.40369752),
    $shortrealtobits(0.3948295),$shortrealtobits(-0.53185457),$shortrealtobits(-0.23099847),$shortrealtobits(-0.13620713),
    $shortrealtobits(0.35436562),$shortrealtobits(-0.4402184),$shortrealtobits(-0.33693582),$shortrealtobits(-0.2595123)
  },
  '{ 
    $shortrealtobits(0.15223147),$shortrealtobits(-0.34290487),$shortrealtobits(-0.030850284),$shortrealtobits(0.13985033),
    $shortrealtobits(-0.2935586),$shortrealtobits(-0.11107563),$shortrealtobits(-0.4647575),$shortrealtobits(-0.2875111),
    $shortrealtobits(0.38672286),$shortrealtobits(0.02345279),$shortrealtobits(-0.40391088),$shortrealtobits(0.0656383),
    $shortrealtobits(0.49548733),$shortrealtobits(-0.55440784),$shortrealtobits(0.033887353),$shortrealtobits(0.32247865),
    $shortrealtobits(-0.0274448),$shortrealtobits(0.5131214),$shortrealtobits(-0.4873458),$shortrealtobits(0.2000358),
    $shortrealtobits(0.23398809),$shortrealtobits(-0.3158826),$shortrealtobits(-0.19164771),$shortrealtobits(0.042201176),
    $shortrealtobits(-0.34807083),$shortrealtobits(0.5057217),$shortrealtobits(-0.2591614),$shortrealtobits(0.38197687),
    $shortrealtobits(0.12573549),$shortrealtobits(0.4112269),$shortrealtobits(0.3208419),$shortrealtobits(-0.17871071),
    $shortrealtobits(-0.18149698),$shortrealtobits(0.106169924),$shortrealtobits(-0.06743195),$shortrealtobits(-0.23321809),
    $shortrealtobits(-0.3164815),$shortrealtobits(-0.32807866),$shortrealtobits(0.41317326),$shortrealtobits(-0.4641507)
  },
  '{ 
    $shortrealtobits(-0.24239427),$shortrealtobits(-0.42859474),$shortrealtobits(0.19741996),$shortrealtobits(0.3538461),
    $shortrealtobits(-0.10305477),$shortrealtobits(-0.22706804),$shortrealtobits(0.05373543),$shortrealtobits(-0.41351315),
    $shortrealtobits(0.096080564),$shortrealtobits(0.43433785),$shortrealtobits(-0.42498827),$shortrealtobits(-0.057621546),
    $shortrealtobits(0.41962942),$shortrealtobits(-0.22363165),$shortrealtobits(-0.44443682),$shortrealtobits(-0.34596953),
    $shortrealtobits(0.21181454),$shortrealtobits(-0.23049511),$shortrealtobits(-0.1405735),$shortrealtobits(-0.048742175),
    $shortrealtobits(0.04695809),$shortrealtobits(0.5682096),$shortrealtobits(-0.14009146),$shortrealtobits(0.46866825),
    $shortrealtobits(0.22046112),$shortrealtobits(0.24097787),$shortrealtobits(0.06242184),$shortrealtobits(0.52168685),
    $shortrealtobits(0.17102224),$shortrealtobits(-0.5925851),$shortrealtobits(0.23579225),$shortrealtobits(-0.046661265),
    $shortrealtobits(-0.19152303),$shortrealtobits(0.3473242),$shortrealtobits(0.054624993),$shortrealtobits(0.05669112),
    $shortrealtobits(0.33725965),$shortrealtobits(0.44505528),$shortrealtobits(-0.3810305),$shortrealtobits(-0.14048809)
  },
  '{ 
    $shortrealtobits(0.490684),$shortrealtobits(-0.25113073),$shortrealtobits(-0.06372514),$shortrealtobits(0.19295976),
    $shortrealtobits(0.25318635),$shortrealtobits(-0.16190057),$shortrealtobits(-0.13138409),$shortrealtobits(0.37241694),
    $shortrealtobits(-0.3673856),$shortrealtobits(0.26368767),$shortrealtobits(-0.016025215),$shortrealtobits(0.16369005),
    $shortrealtobits(0.31231993),$shortrealtobits(-0.4856385),$shortrealtobits(-0.21149161),$shortrealtobits(0.020830657),
    $shortrealtobits(-0.5564368),$shortrealtobits(0.20313919),$shortrealtobits(0.023176435),$shortrealtobits(-0.32155555),
    $shortrealtobits(0.46647778),$shortrealtobits(0.09684472),$shortrealtobits(0.12919457),$shortrealtobits(-0.2421946),
    $shortrealtobits(0.58164805),$shortrealtobits(0.0023954946),$shortrealtobits(0.4012022),$shortrealtobits(0.10600975),
    $shortrealtobits(0.2608932),$shortrealtobits(-0.3185372),$shortrealtobits(0.27170953),$shortrealtobits(-0.15957783),
    $shortrealtobits(-0.053045716),$shortrealtobits(0.4954038),$shortrealtobits(0.00118909),$shortrealtobits(0.24025308),
    $shortrealtobits(-0.04103231),$shortrealtobits(-0.48672074),$shortrealtobits(0.1734871),$shortrealtobits(0.38418496)
  },
  '{ 
    $shortrealtobits(0.15454604),$shortrealtobits(0.17984141),$shortrealtobits(0.44524825),$shortrealtobits(0.043105155),
    $shortrealtobits(-0.18755627),$shortrealtobits(0.021990234),$shortrealtobits(-0.10380355),$shortrealtobits(-0.26898816),
    $shortrealtobits(0.22537687),$shortrealtobits(0.6335219),$shortrealtobits(0.11306679),$shortrealtobits(-0.42392805),
    $shortrealtobits(0.41789424),$shortrealtobits(0.18440373),$shortrealtobits(-0.26662534),$shortrealtobits(-0.059648976),
    $shortrealtobits(-0.29277444),$shortrealtobits(-0.35451117),$shortrealtobits(-0.15591656),$shortrealtobits(0.116857894),
    $shortrealtobits(0.28207308),$shortrealtobits(0.005432398),$shortrealtobits(0.33148432),$shortrealtobits(-0.0070261415),
    $shortrealtobits(0.39463717),$shortrealtobits(-0.32172284),$shortrealtobits(-0.1295887),$shortrealtobits(-0.09193033),
    $shortrealtobits(-0.5661143),$shortrealtobits(-0.03786698),$shortrealtobits(0.76799953),$shortrealtobits(0.06043382),
    $shortrealtobits(0.13988322),$shortrealtobits(0.42010856),$shortrealtobits(0.19835368),$shortrealtobits(0.12132166),
    $shortrealtobits(0.066086106),$shortrealtobits(-0.40939015),$shortrealtobits(0.5085415),$shortrealtobits(-0.16785099)
  },
  '{ 
    $shortrealtobits(0.42606768),$shortrealtobits(-0.0019958187),$shortrealtobits(0.45926684),$shortrealtobits(-0.30377093),
    $shortrealtobits(0.10089745),$shortrealtobits(-0.08821893),$shortrealtobits(-0.069141224),$shortrealtobits(0.097273186),
    $shortrealtobits(0.4593827),$shortrealtobits(0.23145661),$shortrealtobits(-0.19162954),$shortrealtobits(0.16604304),
    $shortrealtobits(-0.38366488),$shortrealtobits(-0.3912803),$shortrealtobits(-0.36000267),$shortrealtobits(0.00020520244),
    $shortrealtobits(-0.23027256),$shortrealtobits(-0.047409166),$shortrealtobits(0.46788874),$shortrealtobits(-0.2827697),
    $shortrealtobits(0.20356654),$shortrealtobits(0.2689787),$shortrealtobits(-0.24982136),$shortrealtobits(-0.5984571),
    $shortrealtobits(0.013728556),$shortrealtobits(-0.38677323),$shortrealtobits(0.7076132),$shortrealtobits(0.063394025),
    $shortrealtobits(0.2181527),$shortrealtobits(0.044587437),$shortrealtobits(-0.24578616),$shortrealtobits(0.019789),
    $shortrealtobits(-0.2932969),$shortrealtobits(-0.24334769),$shortrealtobits(-0.004211317),$shortrealtobits(0.14541727),
    $shortrealtobits(-0.38613987),$shortrealtobits(-0.009719139),$shortrealtobits(-0.054765813),$shortrealtobits(-0.32049784)
  },
  '{ 
    $shortrealtobits(0.08463569),$shortrealtobits(-0.028459765),$shortrealtobits(0.12337867),$shortrealtobits(-0.06956175),
    $shortrealtobits(0.0016338917),$shortrealtobits(0.42841962),$shortrealtobits(-0.12826702),$shortrealtobits(-0.37669548),
    $shortrealtobits(0.29588404),$shortrealtobits(0.11624599),$shortrealtobits(0.084575534),$shortrealtobits(0.11469633),
    $shortrealtobits(-0.16431458),$shortrealtobits(0.19827068),$shortrealtobits(-0.22568557),$shortrealtobits(0.03968863),
    $shortrealtobits(0.13414082),$shortrealtobits(-0.0071593067),$shortrealtobits(-0.38504797),$shortrealtobits(0.059948705),
    $shortrealtobits(-0.040269822),$shortrealtobits(0.40158513),$shortrealtobits(0.124019295),$shortrealtobits(0.18839663),
    $shortrealtobits(0.10122424),$shortrealtobits(-0.22605723),$shortrealtobits(-0.26703632),$shortrealtobits(-0.18116525),
    $shortrealtobits(0.042721126),$shortrealtobits(0.238195),$shortrealtobits(-0.35129508),$shortrealtobits(0.38226596),
    $shortrealtobits(0.079037905),$shortrealtobits(-0.23124313),$shortrealtobits(-0.04188772),$shortrealtobits(-0.22549425),
    $shortrealtobits(0.4201498),$shortrealtobits(0.14541231),$shortrealtobits(-0.5066115),$shortrealtobits(0.11091933)
  },
  '{ 
    $shortrealtobits(-0.033057794),$shortrealtobits(0.1797545),$shortrealtobits(-0.06028022),$shortrealtobits(-0.20314242),
    $shortrealtobits(0.3457859),$shortrealtobits(0.06342284),$shortrealtobits(0.37178937),$shortrealtobits(-0.28544873),
    $shortrealtobits(0.1632409),$shortrealtobits(-0.3149954),$shortrealtobits(-0.1965857),$shortrealtobits(-0.22264002),
    $shortrealtobits(0.3913476),$shortrealtobits(0.103143044),$shortrealtobits(0.017200839),$shortrealtobits(0.043210253),
    $shortrealtobits(-0.098439515),$shortrealtobits(0.43460068),$shortrealtobits(-0.43448249),$shortrealtobits(-0.20542105),
    $shortrealtobits(0.37145624),$shortrealtobits(-0.51306486),$shortrealtobits(-0.44228286),$shortrealtobits(-0.4177145),
    $shortrealtobits(-0.07513606),$shortrealtobits(0.4734206),$shortrealtobits(-0.24991395),$shortrealtobits(-0.28147772),
    $shortrealtobits(0.2472236),$shortrealtobits(0.05909792),$shortrealtobits(-0.26295477),$shortrealtobits(-0.15115547),
    $shortrealtobits(-0.35401952),$shortrealtobits(0.33009097),$shortrealtobits(0.34175363),$shortrealtobits(0.025669228),
    $shortrealtobits(-0.006434837),$shortrealtobits(-0.048552677),$shortrealtobits(-0.4047305),$shortrealtobits(0.6784886)
  },
  '{ 
    $shortrealtobits(0.7937354),$shortrealtobits(-0.49544767),$shortrealtobits(0.024364414),$shortrealtobits(0.2314354),
    $shortrealtobits(0.034607396),$shortrealtobits(-0.24003194),$shortrealtobits(0.1923744),$shortrealtobits(0.16557813),
    $shortrealtobits(0.13640246),$shortrealtobits(0.35691404),$shortrealtobits(0.16527343),$shortrealtobits(-0.34459984),
    $shortrealtobits(-0.37019402),$shortrealtobits(0.43146193),$shortrealtobits(-0.20775588),$shortrealtobits(0.01262055),
    $shortrealtobits(-0.3677737),$shortrealtobits(-0.5966505),$shortrealtobits(-0.29081666),$shortrealtobits(0.13032885),
    $shortrealtobits(0.20107013),$shortrealtobits(0.17280626),$shortrealtobits(0.49653068),$shortrealtobits(-0.15279295),
    $shortrealtobits(0.033706814),$shortrealtobits(-0.3438691),$shortrealtobits(-0.78677404),$shortrealtobits(-0.02825357),
    $shortrealtobits(-0.5479744),$shortrealtobits(-0.45100507),$shortrealtobits(-0.43634033),$shortrealtobits(-0.11329835),
    $shortrealtobits(-0.31753203),$shortrealtobits(0.15156679),$shortrealtobits(-0.039174255),$shortrealtobits(0.046175264),
    $shortrealtobits(0.13501824),$shortrealtobits(-0.5412288),$shortrealtobits(-0.010190201),$shortrealtobits(-0.29624826)
  },
  '{ 
    $shortrealtobits(0.5606924),$shortrealtobits(-0.48780832),$shortrealtobits(-0.6902587),$shortrealtobits(-0.05174905),
    $shortrealtobits(0.013552625),$shortrealtobits(0.5909365),$shortrealtobits(0.10735167),$shortrealtobits(0.40221697),
    $shortrealtobits(0.86055726),$shortrealtobits(0.3002334),$shortrealtobits(-0.50604147),$shortrealtobits(0.04779879),
    $shortrealtobits(-0.060957156),$shortrealtobits(-0.07422514),$shortrealtobits(0.14914711),$shortrealtobits(0.47260165),
    $shortrealtobits(0.27691835),$shortrealtobits(0.22121453),$shortrealtobits(-0.17155771),$shortrealtobits(-0.3193869),
    $shortrealtobits(-0.34348857),$shortrealtobits(0.32767367),$shortrealtobits(-0.3960305),$shortrealtobits(-0.6109),
    $shortrealtobits(0.19084723),$shortrealtobits(-0.26179007),$shortrealtobits(-0.24973789),$shortrealtobits(0.24757363),
    $shortrealtobits(-0.28460997),$shortrealtobits(0.036036473),$shortrealtobits(-0.4214159),$shortrealtobits(-0.23020749),
    $shortrealtobits(0.5647155),$shortrealtobits(-0.3486379),$shortrealtobits(-0.53194076),$shortrealtobits(-0.31539616),
    $shortrealtobits(-0.2743365),$shortrealtobits(-0.39277902),$shortrealtobits(-0.5917949),$shortrealtobits(-0.22401291)
  },
  '{ 
    $shortrealtobits(-0.03746161),$shortrealtobits(0.015650779),$shortrealtobits(0.16271508),$shortrealtobits(-0.40732065),
    $shortrealtobits(-0.4687111),$shortrealtobits(-0.19836037),$shortrealtobits(0.22099137),$shortrealtobits(0.0342536),
    $shortrealtobits(-0.15580644),$shortrealtobits(0.12315232),$shortrealtobits(0.11206117),$shortrealtobits(0.25329062),
    $shortrealtobits(-0.1777647),$shortrealtobits(0.41931522),$shortrealtobits(-0.33521277),$shortrealtobits(-0.031493574),
    $shortrealtobits(0.13866709),$shortrealtobits(-0.3518911),$shortrealtobits(-0.56424546),$shortrealtobits(0.08449142),
    $shortrealtobits(-0.35041562),$shortrealtobits(-0.020378472),$shortrealtobits(-0.5165471),$shortrealtobits(-0.29305384),
    $shortrealtobits(-0.44812426),$shortrealtobits(0.33359134),$shortrealtobits(0.16313045),$shortrealtobits(-0.20164873),
    $shortrealtobits(-0.137697),$shortrealtobits(0.41990793),$shortrealtobits(0.13508089),$shortrealtobits(0.009772274),
    $shortrealtobits(-0.2617505),$shortrealtobits(-0.30223948),$shortrealtobits(-0.10970777),$shortrealtobits(-0.46040145),
    $shortrealtobits(-0.3317712),$shortrealtobits(-0.45670828),$shortrealtobits(-0.41823596),$shortrealtobits(0.29807115)
  },
  '{ 
    $shortrealtobits(0.2831055),$shortrealtobits(-0.029303966),$shortrealtobits(-0.6298296),$shortrealtobits(-0.102993116),
    $shortrealtobits(0.43879044),$shortrealtobits(0.5057988),$shortrealtobits(0.1215451),$shortrealtobits(0.33902916),
    $shortrealtobits(0.88066554),$shortrealtobits(0.4748264),$shortrealtobits(-0.6082616),$shortrealtobits(-0.21927457),
    $shortrealtobits(-0.4199076),$shortrealtobits(-0.4753914),$shortrealtobits(0.11814689),$shortrealtobits(0.06205031),
    $shortrealtobits(0.21575926),$shortrealtobits(-0.5039627),$shortrealtobits(0.010370975),$shortrealtobits(0.09787602),
    $shortrealtobits(-0.029063934),$shortrealtobits(0.12573943),$shortrealtobits(-0.13483576),$shortrealtobits(-0.33243716),
    $shortrealtobits(-0.0036280924),$shortrealtobits(-0.3922925),$shortrealtobits(-0.2850565),$shortrealtobits(0.0071651377),
    $shortrealtobits(-0.5975193),$shortrealtobits(-0.2840353),$shortrealtobits(-0.5521324),$shortrealtobits(0.40599948),
    $shortrealtobits(-0.14195292),$shortrealtobits(0.21745202),$shortrealtobits(-1.0599755),$shortrealtobits(-0.2405033),
    $shortrealtobits(-0.12961465),$shortrealtobits(-0.61987245),$shortrealtobits(0.23306897),$shortrealtobits(-0.3851709)
	}
};

    accel_dot #(
        .ROWS(ROWS),
        .COLS(COLS)
    ) accel_dot0 (
    
		// AXI4-Stream Interface
		.clk(clk),
		.rst(rst),
		
        .weights(weights),

        .INPUT_AXIS_TDATA(INPUT_AXIS_TDATA),
        .INPUT_AXIS_TLAST(INPUT_AXIS_TLAST),
        .INPUT_AXIS_TVALID(INPUT_AXIS_TVALID),
        .INPUT_AXIS_TREADY(INPUT_AXIS_TREADY),
                            
        .OUTPUT_AXIS_TDATA(OUTPUT_AXIS_TDATA),
        .OUTPUT_AXIS_TLAST(OUTPUT_AXIS_TLAST),
        .OUTPUT_AXIS_TVALID(OUTPUT_AXIS_TVALID),
        .OUTPUT_AXIS_TREADY(OUTPUT_AXIS_TREADY) 	

    );

    
endmodule
